/******************************************************************************

   The MIT License (MIT)

   Copyright (c) 2015 Embedded Micro

   Permission is hereby granted, free of charge, to any person obtaining a copy
   of this software and associated documentation files (the "Software"), to deal
   in the Software without restriction, including without limitation the rights
   to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
   copies of the Software, and to permit persons to whom the Software is
   furnished to do so, subject to the following conditions:

   The above copyright notice and this permission notice shall be included in
   all copies or substantial portions of the Software.

   THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
   IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
   FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
   AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
   LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
   OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
   THE SOFTWARE.

   *****************************************************************************

   This module is a simple single port RAM. This RAM is implemented in such a
   way that Xilinx's tools will recognize it as a RAM and implement large
   instances in block RAM instead of flip-flops.
   
   The parameter SIZE is used to specify the word size. That is the size of 
   each entry in the RAM.
   
   The parameter DEPTH is used to specify how many entries are in the RAM.
   
   read_data outputs the value of the entry pointed to by address in the previous
   clock cycle. That means to read address 10, you would set address to be 10
   and wait one cycle for its value to show up. The RAM is always reading whatever
   address is. If you don't need to read, just ignore this value.
   
   To write, set write_en to 1, write_data to the value to write,
   and address to the address you want to write.
   
   If you read and write the same address, the first clock cycle the address will
   be written, the second clock cycle the old value will be output on read_data,
   and on the third clock cycle the newly updated value will be output on 
   read_data.
*/

module simple_ram #(
    parameter SIZE = 8,  // size of each entry
    parameter DEPTH = 80,  // number of entries
    parameter MEM_INIT_FILE = 0
  )(
    input clk,                         // clock
    input [$clog2(DEPTH)-1:0] address, // address to read or write
    output reg [SIZE-1:0] read_data,   // data read
    input [SIZE-1:0] write_data,       // data to write
    input write_en                     // write enable (1 = write)
  );
  
  reg [SIZE-1:0] ram [DEPTH-1:0];      // memory array
  
initial begin
  //if (MEM_INIT_FILE != "") begin
   // $readmemb("MEM_INT_FILE", ram);
  //end
  
case(MEM_INIT_FILE)

0 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "n";
ram[5] = "e";
ram[6] = "i";
ram[7] = "g";
ram[8] = "h";
ram[9] = "b";
ram[10] = "o";
ram[11] = "u";
ram[12] = "r";
ram[13] = "i";
ram[14] = "n";
ram[15] = "g";
ram[16] = " ";
ram[17] = "k";
ram[18] = "i";
ram[19] = "n";
ram[20] = "g";
ram[21] = "d";
ram[22] = "o";
ram[23] = "m";
ram[24] = " ";
ram[25] = "h";
ram[26] = "a";
ram[27] = "s";
ram[28] = " ";
ram[29] = "b";
ram[30] = "e";
ram[31] = "e";
ram[32] = "n";
ram[33] = " ";
ram[34] = "w";
ram[35] = "e";
ram[36] = "a";
ram[37] = "k";
ram[38] = "e";
ram[39] = "n";
ram[40] = "e";
ram[41] = "d";
ram[42] = ".";
ram[43] = " ";
ram[44] = "I";
ram[45] = "n";
ram[46] = "v";
ram[47] = "a";
ram[48] = "d";
ram[49] = "e";
ram[50] = " ";
ram[51] = "t";
ram[52] = "h";
ram[53] = "e";
ram[54] = " ";
ram[55] = "n";
ram[56] = "e";
ram[57] = "i";
ram[58] = "g";
ram[59] = "h";
ram[60] = "b";
ram[61] = "o";
ram[62] = "u";
ram[63] = "r";
ram[64] = "i";
ram[65] = "n";
ram[66] = "g";
ram[67] = " ";
ram[68] = "k";
ram[69] = "i";
ram[70] = "n";
ram[71] = "g";
ram[72] = "d";
ram[73] = "o";
ram[74] = "m";
ram[75] = "?";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
1 : begin
ram[0] = "Y";
ram[1] = "o";
ram[2] = "u";
ram[3] = "r";
ram[4] = " ";
ram[5] = "m";
ram[6] = "i";
ram[7] = "l";
ram[8] = "i";
ram[9] = "t";
ram[10] = "a";
ram[11] = "r";
ram[12] = "y";
ram[13] = " ";
ram[14] = "w";
ram[15] = "i";
ram[16] = "s";
ram[17] = "h";
ram[18] = "e";
ram[19] = "s";
ram[20] = " ";
ram[21] = "t";
ram[22] = "o";
ram[23] = " ";
ram[24] = "c";
ram[25] = "o";
ram[26] = "n";
ram[27] = "d";
ram[28] = "u";
ram[29] = "c";
ram[30] = "t";
ram[31] = " ";
ram[32] = "a";
ram[33] = " ";
ram[34] = "h";
ram[35] = "u";
ram[36] = "n";
ram[37] = "t";
ram[38] = " ";
ram[39] = "i";
ram[40] = "n";
ram[41] = " ";
ram[42] = "t";
ram[43] = "h";
ram[44] = "e";
ram[45] = " ";
ram[46] = "w";
ram[47] = "o";
ram[48] = "o";
ram[49] = "d";
ram[50] = "s";
ram[51] = ".";
ram[52] = " ";
ram[53] = "J";
ram[54] = "o";
ram[55] = "i";
ram[56] = "n";
ram[57] = " ";
ram[58] = "t";
ram[59] = "h";
ram[60] = "e";
ram[61] = "m";
ram[62] = "?";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
2 : begin
ram[0] = "Y";
ram[1] = "o";
ram[2] = "u";
ram[3] = "r";
ram[4] = " ";
ram[5] = "e";
ram[6] = "n";
ram[7] = "e";
ram[8] = "m";
ram[9] = "i";
ram[10] = "e";
ram[11] = "s";
ram[12] = " ";
ram[13] = "w";
ram[14] = "a";
ram[15] = "n";
ram[16] = "t";
ram[17] = " ";
ram[18] = "t";
ram[19] = "o";
ram[20] = " ";
ram[21] = "s";
ram[22] = "i";
ram[23] = "g";
ram[24] = "n";
ram[25] = " ";
ram[26] = "a";
ram[27] = " ";
ram[28] = "p";
ram[29] = "e";
ram[30] = "a";
ram[31] = "c";
ram[32] = "e";
ram[33] = " ";
ram[34] = "t";
ram[35] = "r";
ram[36] = "e";
ram[37] = "a";
ram[38] = "t";
ram[39] = "y";
ram[40] = " ";
ram[41] = "t";
ram[42] = "o";
ram[43] = " ";
ram[44] = "p";
ram[45] = "r";
ram[46] = "e";
ram[47] = "v";
ram[48] = "e";
ram[49] = "n";
ram[50] = "t";
ram[51] = " ";
ram[52] = "w";
ram[53] = "a";
ram[54] = "r";
ram[55] = ".";
ram[56] = " ";
ram[57] = "S";
ram[58] = "i";
ram[59] = "g";
ram[60] = "n";
ram[61] = " ";
ram[62] = "t";
ram[63] = "h";
ram[64] = "e";
ram[65] = " ";
ram[66] = "t";
ram[67] = "r";
ram[68] = "e";
ram[69] = "a";
ram[70] = "t";
ram[71] = "y";
ram[72] = "?";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
3 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "c";
ram[5] = "h";
ram[6] = "u";
ram[7] = "r";
ram[8] = "c";
ram[9] = "h";
ram[10] = " ";
ram[11] = "w";
ram[12] = "a";
ram[13] = "n";
ram[14] = "t";
ram[15] = "s";
ram[16] = " ";
ram[17] = "t";
ram[18] = "o";
ram[19] = " ";
ram[20] = "s";
ram[21] = "t";
ram[22] = "a";
ram[23] = "r";
ram[24] = "t";
ram[25] = " ";
ram[26] = "a";
ram[27] = " ";
ram[28] = "w";
ram[29] = "a";
ram[30] = "r";
ram[31] = " ";
ram[32] = "w";
ram[33] = "i";
ram[34] = "t";
ram[35] = "h";
ram[36] = " ";
ram[37] = "t";
ram[38] = "h";
ram[39] = "e";
ram[40] = " ";
ram[41] = "p";
ram[42] = "a";
ram[43] = "g";
ram[44] = "a";
ram[45] = "n";
ram[46] = "s";
ram[47] = ",";
ram[48] = " ";
ram[49] = "l";
ram[50] = "e";
ram[51] = "t";
ram[52] = " ";
ram[53] = "t";
ram[54] = "h";
ram[55] = "e";
ram[56] = "m";
ram[57] = "?";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
4 : begin
ram[0] = "S";
ram[1] = "i";
ram[2] = "r";
ram[3] = "e";
ram[4] = ",";
ram[5] = " ";
ram[6] = "o";
ram[7] = "u";
ram[8] = "r";
ram[9] = " ";
ram[10] = "m";
ram[11] = "e";
ram[12] = "n";
ram[13] = " ";
ram[14] = "g";
ram[15] = "r";
ram[16] = "o";
ram[17] = "w";
ram[18] = " ";
ram[19] = "r";
ram[20] = "e";
ram[21] = "s";
ram[22] = "t";
ram[23] = "l";
ram[24] = "e";
ram[25] = "s";
ram[26] = "s";
ram[27] = ".";
ram[28] = " ";
ram[29] = "S";
ram[30] = "h";
ram[31] = "a";
ram[32] = "l";
ram[33] = "l";
ram[34] = " ";
ram[35] = "w";
ram[36] = "e";
ram[37] = " ";
ram[38] = "t";
ram[39] = "u";
ram[40] = "r";
ram[41] = "n";
ram[42] = " ";
ram[43] = "t";
ram[44] = "h";
ram[45] = "e";
ram[46] = "i";
ram[47] = "r";
ram[48] = " ";
ram[49] = "w";
ram[50] = "a";
ram[51] = "t";
ram[52] = "e";
ram[53] = "r";
ram[54] = " ";
ram[55] = "i";
ram[56] = "n";
ram[57] = "t";
ram[58] = "o";
ram[59] = " ";
ram[60] = "w";
ram[61] = "i";
ram[62] = "n";
ram[63] = "e";
ram[64] = "?";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
5 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "c";
ram[5] = "h";
ram[6] = "u";
ram[7] = "r";
ram[8] = "c";
ram[9] = "h";
ram[10] = " ";
ram[11] = "i";
ram[12] = "s";
ram[13] = " ";
ram[14] = "l";
ram[15] = "a";
ram[16] = "c";
ram[17] = "k";
ram[18] = "i";
ram[19] = "n";
ram[20] = "g";
ram[21] = " ";
ram[22] = "m";
ram[23] = "a";
ram[24] = "n";
ram[25] = "p";
ram[26] = "o";
ram[27] = "w";
ram[28] = "e";
ram[29] = "r";
ram[30] = ".";
ram[31] = " ";
ram[32] = "R";
ram[33] = "e";
ram[34] = "c";
ram[35] = "r";
ram[36] = "u";
ram[37] = "i";
ram[38] = "t";
ram[39] = " ";
ram[40] = "m";
ram[41] = "o";
ram[42] = "r";
ram[43] = "e";
ram[44] = " ";
ram[45] = "c";
ram[46] = "h";
ram[47] = "u";
ram[48] = "r";
ram[49] = "c";
ram[50] = "h";
ram[51] = " ";
ram[52] = "o";
ram[53] = "f";
ram[54] = "f";
ram[55] = "i";
ram[56] = "c";
ram[57] = "i";
ram[58] = "a";
ram[59] = "l";
ram[60] = "s";
ram[61] = " ";
ram[62] = "f";
ram[63] = "r";
ram[64] = "o";
ram[65] = "m";
ram[66] = " ";
ram[67] = "t";
ram[68] = "h";
ram[69] = "e";
ram[70] = " ";
ram[71] = "p";
ram[72] = "e";
ram[73] = "o";
ram[74] = "p";
ram[75] = "l";
ram[76] = "e";
ram[77] = "?";
ram[78] = " ";
ram[79] = " ";
end
6 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "c";
ram[5] = "h";
ram[6] = "u";
ram[7] = "r";
ram[8] = "c";
ram[9] = "h";
ram[10] = " ";
ram[11] = "w";
ram[12] = "o";
ram[13] = "u";
ram[14] = "l";
ram[15] = "d";
ram[16] = " ";
ram[17] = "l";
ram[18] = "i";
ram[19] = "k";
ram[20] = "e";
ram[21] = " ";
ram[22] = "t";
ram[23] = "o";
ram[24] = " ";
ram[25] = "b";
ram[26] = "u";
ram[27] = "i";
ram[28] = "l";
ram[29] = "d";
ram[30] = " ";
ram[31] = "s";
ram[32] = "c";
ram[33] = "h";
ram[34] = "o";
ram[35] = "o";
ram[36] = "l";
ram[37] = "s";
ram[38] = " ";
ram[39] = "f";
ram[40] = "o";
ram[41] = "r";
ram[42] = " ";
ram[43] = "t";
ram[44] = "h";
ram[45] = "e";
ram[46] = " ";
ram[47] = "p";
ram[48] = "e";
ram[49] = "o";
ram[50] = "p";
ram[51] = "l";
ram[52] = "e";
ram[53] = ".";
ram[54] = " ";
ram[55] = "A";
ram[56] = "l";
ram[57] = "l";
ram[58] = "o";
ram[59] = "w";
ram[60] = " ";
ram[61] = "t";
ram[62] = "h";
ram[63] = "e";
ram[64] = "m";
ram[65] = "?";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
7 : begin
ram[0] = "A";
ram[1] = " ";
ram[2] = "f";
ram[3] = "e";
ram[4] = "w";
ram[5] = " ";
ram[6] = "m";
ram[7] = "o";
ram[8] = "n";
ram[9] = "k";
ram[10] = "s";
ram[11] = " ";
ram[12] = "h";
ram[13] = "a";
ram[14] = "v";
ram[15] = "e";
ram[16] = " ";
ram[17] = "b";
ram[18] = "e";
ram[19] = "e";
ram[20] = "n";
ram[21] = " ";
ram[22] = "f";
ram[23] = "o";
ram[24] = "u";
ram[25] = "n";
ram[26] = "d";
ram[27] = " ";
ram[28] = "b";
ram[29] = "e";
ram[30] = "h";
ram[31] = "a";
ram[32] = "v";
ram[33] = "i";
ram[34] = "n";
ram[35] = "g";
ram[36] = " ";
ram[37] = "l";
ram[38] = "i";
ram[39] = "k";
ram[40] = "e";
ram[41] = " ";
ram[42] = "d";
ram[43] = "u";
ram[44] = "c";
ram[45] = "k";
ram[46] = "s";
ram[47] = " ";
ram[48] = "i";
ram[49] = "n";
ram[50] = " ";
ram[51] = "t";
ram[52] = "h";
ram[53] = "e";
ram[54] = " ";
ram[55] = "s";
ram[56] = "q";
ram[57] = "u";
ram[58] = "a";
ram[59] = "r";
ram[60] = "e";
ram[61] = ",";
ram[62] = " ";
ram[63] = "l";
ram[64] = "o";
ram[65] = "c";
ram[66] = "k";
ram[67] = " ";
ram[68] = "t";
ram[69] = "h";
ram[70] = "e";
ram[71] = "m";
ram[72] = " ";
ram[73] = "u";
ram[74] = "p";
ram[75] = "?";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
8 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "p";
ram[5] = "o";
ram[6] = "p";
ram[7] = "e";
ram[8] = " ";
ram[9] = "r";
ram[10] = "e";
ram[11] = "q";
ram[12] = "u";
ram[13] = "e";
ram[14] = "s";
ram[15] = "t";
ram[16] = "s";
ram[17] = " ";
ram[18] = "t";
ram[19] = "o";
ram[20] = " ";
ram[21] = "d";
ram[22] = "e";
ram[23] = "c";
ram[24] = "l";
ram[25] = "a";
ram[26] = "r";
ram[27] = "e";
ram[28] = " ";
ram[29] = "2";
ram[30] = "5";
ram[31] = "t";
ram[32] = "h";
ram[33] = " ";
ram[34] = "D";
ram[35] = "e";
ram[36] = "c";
ram[37] = "e";
ram[38] = "m";
ram[39] = "b";
ram[40] = "e";
ram[41] = "r";
ram[42] = " ";
ram[43] = "a";
ram[44] = " ";
ram[45] = "n";
ram[46] = "e";
ram[47] = "w";
ram[48] = " ";
ram[49] = "h";
ram[50] = "o";
ram[51] = "l";
ram[52] = "i";
ram[53] = "d";
ram[54] = "a";
ram[55] = "y";
ram[56] = ",";
ram[57] = " ";
ram[58] = "C";
ram[59] = "h";
ram[60] = "r";
ram[61] = "i";
ram[62] = "s";
ram[63] = "t";
ram[64] = " ";
ram[65] = "M";
ram[66] = "a";
ram[67] = "s";
ram[68] = "s";
ram[69] = ".";
ram[70] = " ";
ram[71] = "A";
ram[72] = "g";
ram[73] = "r";
ram[74] = "e";
ram[75] = "e";
ram[76] = "?";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
9 : begin
ram[0] = "I";
ram[1] = "s";
ram[2] = " ";
ram[3] = "t";
ram[4] = "h";
ram[5] = "e";
ram[6] = " ";
ram[7] = "e";
ram[8] = "a";
ram[9] = "r";
ram[10] = "t";
ram[11] = "h";
ram[12] = " ";
ram[13] = "r";
ram[14] = "o";
ram[15] = "u";
ram[16] = "n";
ram[17] = "d";
ram[18] = "?";
ram[19] = " ";
ram[20] = " ";
ram[21] = " ";
ram[22] = " ";
ram[23] = " ";
ram[24] = " ";
ram[25] = " ";
ram[26] = " ";
ram[27] = " ";
ram[28] = " ";
ram[29] = " ";
ram[30] = " ";
ram[31] = " ";
ram[32] = " ";
ram[33] = " ";
ram[34] = " ";
ram[35] = " ";
ram[36] = " ";
ram[37] = " ";
ram[38] = " ";
ram[39] = " ";
ram[40] = " ";
ram[41] = " ";
ram[42] = " ";
ram[43] = " ";
ram[44] = " ";
ram[45] = " ";
ram[46] = " ";
ram[47] = " ";
ram[48] = " ";
ram[49] = " ";
ram[50] = " ";
ram[51] = " ";
ram[52] = " ";
ram[53] = " ";
ram[54] = " ";
ram[55] = " ";
ram[56] = " ";
ram[57] = " ";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
10 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "p";
ram[5] = "e";
ram[6] = "o";
ram[7] = "p";
ram[8] = "l";
ram[9] = "e";
ram[10] = " ";
ram[11] = "a";
ram[12] = "r";
ram[13] = "e";
ram[14] = " ";
ram[15] = "l";
ram[16] = "o";
ram[17] = "s";
ram[18] = "i";
ram[19] = "n";
ram[20] = "g";
ram[21] = " ";
ram[22] = "f";
ram[23] = "a";
ram[24] = "i";
ram[25] = "t";
ram[26] = "h";
ram[27] = " ";
ram[28] = "i";
ram[29] = "n";
ram[30] = " ";
ram[31] = "t";
ram[32] = "h";
ram[33] = "e";
ram[34] = " ";
ram[35] = "c";
ram[36] = "h";
ram[37] = "u";
ram[38] = "r";
ram[39] = "c";
ram[40] = "h";
ram[41] = ".";
ram[42] = " ";
ram[43] = "E";
ram[44] = "s";
ram[45] = "t";
ram[46] = "a";
ram[47] = "b";
ram[48] = "l";
ram[49] = "i";
ram[50] = "s";
ram[51] = "h";
ram[52] = " ";
ram[53] = "m";
ram[54] = "o";
ram[55] = "r";
ram[56] = "e";
ram[57] = " ";
ram[58] = "c";
ram[59] = "h";
ram[60] = "u";
ram[61] = "r";
ram[62] = "c";
ram[63] = "h";
ram[64] = "e";
ram[65] = "s";
ram[66] = "?";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
11 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "p";
ram[5] = "r";
ram[6] = "i";
ram[7] = "e";
ram[8] = "s";
ram[9] = "t";
ram[10] = "s";
ram[11] = " ";
ram[12] = "r";
ram[13] = "e";
ram[14] = "q";
ram[15] = "u";
ram[16] = "i";
ram[17] = "r";
ram[18] = "e";
ram[19] = " ";
ram[20] = "m";
ram[21] = "o";
ram[22] = "r";
ram[23] = "e";
ram[24] = " ";
ram[25] = "f";
ram[26] = "u";
ram[27] = "n";
ram[28] = "d";
ram[29] = "s";
ram[30] = " ";
ram[31] = "t";
ram[32] = "o";
ram[33] = " ";
ram[34] = "m";
ram[35] = "a";
ram[36] = "i";
ram[37] = "n";
ram[38] = "t";
ram[39] = "a";
ram[40] = "i";
ram[41] = "n";
ram[42] = " ";
ram[43] = "t";
ram[44] = "h";
ram[45] = "e";
ram[46] = "i";
ram[47] = "r";
ram[48] = " ";
ram[49] = "l";
ram[50] = "i";
ram[51] = "f";
ram[52] = "e";
ram[53] = "s";
ram[54] = "t";
ram[55] = "y";
ram[56] = "l";
ram[57] = "e";
ram[58] = "s";
ram[59] = ".";
ram[60] = " ";
ram[61] = "D";
ram[62] = "o";
ram[63] = "n";
ram[64] = "a";
ram[65] = "t";
ram[66] = "e";
ram[67] = " ";
ram[68] = "t";
ram[69] = "o";
ram[70] = " ";
ram[71] = "t";
ram[72] = "h";
ram[73] = "e";
ram[74] = "m";
ram[75] = "?";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
12 : begin
ram[0] = "Y";
ram[1] = "o";
ram[2] = "u";
ram[3] = "r";
ram[4] = " ";
ram[5] = "a";
ram[6] = "d";
ram[7] = "v";
ram[8] = "i";
ram[9] = "s";
ram[10] = "o";
ram[11] = "r";
ram[12] = "s";
ram[13] = " ";
ram[14] = "r";
ram[15] = "e";
ram[16] = "c";
ram[17] = "o";
ram[18] = "m";
ram[19] = "m";
ram[20] = "e";
ram[21] = "n";
ram[22] = "d";
ram[23] = " ";
ram[24] = "y";
ram[25] = "o";
ram[26] = "u";
ram[27] = " ";
ram[28] = "i";
ram[29] = "n";
ram[30] = "v";
ram[31] = "e";
ram[32] = "s";
ram[33] = "t";
ram[34] = " ";
ram[35] = "i";
ram[36] = "n";
ram[37] = " ";
ram[38] = "g";
ram[39] = "o";
ram[40] = "l";
ram[41] = "d";
ram[42] = " ";
ram[43] = "i";
ram[44] = "n";
ram[45] = "s";
ram[46] = "t";
ram[47] = "e";
ram[48] = "a";
ram[49] = "d";
ram[50] = " ";
ram[51] = "o";
ram[52] = "f";
ram[53] = " ";
ram[54] = "t";
ram[55] = "h";
ram[56] = "e";
ram[57] = " ";
ram[58] = "c";
ram[59] = "h";
ram[60] = "u";
ram[61] = "r";
ram[62] = "c";
ram[63] = "h";
ram[64] = ".";
ram[65] = " ";
ram[66] = "I";
ram[67] = "n";
ram[68] = "v";
ram[69] = "e";
ram[70] = "s";
ram[71] = "t";
ram[72] = "?";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
13 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "c";
ram[5] = "h";
ram[6] = "u";
ram[7] = "r";
ram[8] = "c";
ram[9] = "h";
ram[10] = " ";
ram[11] = "w";
ram[12] = "a";
ram[13] = "n";
ram[14] = "t";
ram[15] = "s";
ram[16] = " ";
ram[17] = "t";
ram[18] = "o";
ram[19] = " ";
ram[20] = "i";
ram[21] = "m";
ram[22] = "p";
ram[23] = "o";
ram[24] = "s";
ram[25] = "e";
ram[26] = " ";
ram[27] = "m";
ram[28] = "a";
ram[29] = "n";
ram[30] = "d";
ram[31] = "a";
ram[32] = "t";
ram[33] = "o";
ram[34] = "r";
ram[35] = "y";
ram[36] = " ";
ram[37] = "d";
ram[38] = "o";
ram[39] = "n";
ram[40] = "a";
ram[41] = "t";
ram[42] = "i";
ram[43] = "o";
ram[44] = "n";
ram[45] = "s";
ram[46] = ",";
ram[47] = " ";
ram[48] = "y";
ram[49] = "a";
ram[50] = "y";
ram[51] = " ";
ram[52] = "o";
ram[53] = "r";
ram[54] = " ";
ram[55] = "n";
ram[56] = "a";
ram[57] = "y";
ram[58] = "?";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
14 : begin
ram[0] = "W";
ram[1] = "e";
ram[2] = " ";
ram[3] = "m";
ram[4] = "u";
ram[5] = "s";
ram[6] = "t";
ram[7] = " ";
ram[8] = "i";
ram[9] = "n";
ram[10] = "c";
ram[11] = "r";
ram[12] = "e";
ram[13] = "a";
ram[14] = "s";
ram[15] = "e";
ram[16] = " ";
ram[17] = "o";
ram[18] = "u";
ram[19] = "r";
ram[20] = " ";
ram[21] = "m";
ram[22] = "i";
ram[23] = "l";
ram[24] = "i";
ram[25] = "t";
ram[26] = "a";
ram[27] = "r";
ram[28] = "y";
ram[29] = " ";
ram[30] = "m";
ram[31] = "i";
ram[32] = "g";
ram[33] = "h";
ram[34] = "t";
ram[35] = ".";
ram[36] = " ";
ram[37] = "E";
ram[38] = "n";
ram[39] = "l";
ram[40] = "i";
ram[41] = "s";
ram[42] = "t";
ram[43] = " ";
ram[44] = "c";
ram[45] = "h";
ram[46] = "i";
ram[47] = "l";
ram[48] = "d";
ram[49] = "r";
ram[50] = "e";
ram[51] = "n";
ram[52] = "?";
ram[53] = " ";
ram[54] = " ";
ram[55] = " ";
ram[56] = " ";
ram[57] = " ";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
15 : begin
ram[0] = "W";
ram[1] = "e";
ram[2] = " ";
ram[3] = "n";
ram[4] = "e";
ram[5] = "e";
ram[6] = "d";
ram[7] = " ";
ram[8] = "m";
ram[9] = "o";
ram[10] = "r";
ram[11] = "e";
ram[12] = " ";
ram[13] = "s";
ram[14] = "o";
ram[15] = "l";
ram[16] = "d";
ram[17] = "i";
ram[18] = "e";
ram[19] = "r";
ram[20] = "s";
ram[21] = ".";
ram[22] = " ";
ram[23] = "R";
ram[24] = "e";
ram[25] = "c";
ram[26] = "r";
ram[27] = "u";
ram[28] = "i";
ram[29] = "t";
ram[30] = " ";
ram[31] = "t";
ram[32] = "h";
ram[33] = "e";
ram[34] = " ";
ram[35] = "w";
ram[36] = "o";
ram[37] = "m";
ram[38] = "e";
ram[39] = "n";
ram[40] = "?";
ram[41] = " ";
ram[42] = " ";
ram[43] = " ";
ram[44] = " ";
ram[45] = " ";
ram[46] = " ";
ram[47] = " ";
ram[48] = " ";
ram[49] = " ";
ram[50] = " ";
ram[51] = " ";
ram[52] = " ";
ram[53] = " ";
ram[54] = " ";
ram[55] = " ";
ram[56] = " ";
ram[57] = " ";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
16 : begin
ram[0] = "Y";
ram[1] = "o";
ram[2] = "u";
ram[3] = "r";
ram[4] = " ";
ram[5] = "g";
ram[6] = "e";
ram[7] = "n";
ram[8] = "e";
ram[9] = "r";
ram[10] = "a";
ram[11] = "l";
ram[12] = " ";
ram[13] = "h";
ram[14] = "a";
ram[15] = "s";
ram[16] = " ";
ram[17] = "b";
ram[18] = "e";
ram[19] = "e";
ram[20] = "n";
ram[21] = " ";
ram[22] = "c";
ram[23] = "h";
ram[24] = "a";
ram[25] = "l";
ram[26] = "l";
ram[27] = "e";
ram[28] = "n";
ram[29] = "g";
ram[30] = "e";
ram[31] = "d";
ram[32] = " ";
ram[33] = "t";
ram[34] = "o";
ram[35] = " ";
ram[36] = "a";
ram[37] = " ";
ram[38] = "d";
ram[39] = "u";
ram[40] = "e";
ram[41] = "l";
ram[42] = ".";
ram[43] = " ";
ram[44] = "A";
ram[45] = "l";
ram[46] = "l";
ram[47] = "o";
ram[48] = "w";
ram[49] = " ";
ram[50] = "h";
ram[51] = "i";
ram[52] = "m";
ram[53] = " ";
ram[54] = "t";
ram[55] = "o";
ram[56] = " ";
ram[57] = "t";
ram[58] = "a";
ram[59] = "k";
ram[60] = "e";
ram[61] = " ";
ram[62] = "u";
ram[63] = "p";
ram[64] = " ";
ram[65] = "t";
ram[66] = "h";
ram[67] = "e";
ram[68] = " ";
ram[69] = "d";
ram[70] = "u";
ram[71] = "e";
ram[72] = "l";
ram[73] = "?";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
17 : begin
ram[0] = "Y";
ram[1] = "o";
ram[2] = "u";
ram[3] = "r";
ram[4] = " ";
ram[5] = "s";
ram[6] = "o";
ram[7] = "l";
ram[8] = "d";
ram[9] = "i";
ram[10] = "e";
ram[11] = "r";
ram[12] = "s";
ram[13] = " ";
ram[14] = "h";
ram[15] = "a";
ram[16] = "v";
ram[17] = "e";
ram[18] = " ";
ram[19] = "b";
ram[20] = "e";
ram[21] = "e";
ram[22] = "n";
ram[23] = " ";
ram[24] = "f";
ram[25] = "o";
ram[26] = "u";
ram[27] = "n";
ram[28] = "d";
ram[29] = " ";
ram[30] = "r";
ram[31] = "a";
ram[32] = "p";
ram[33] = "i";
ram[34] = "n";
ram[35] = "g";
ram[36] = " ";
ram[37] = "w";
ram[38] = "o";
ram[39] = "m";
ram[40] = "e";
ram[41] = "n";
ram[42] = ".";
ram[43] = " ";
ram[44] = "E";
ram[45] = "x";
ram[46] = "e";
ram[47] = "c";
ram[48] = "u";
ram[49] = "t";
ram[50] = "e";
ram[51] = " ";
ram[52] = "t";
ram[53] = "h";
ram[54] = "e";
ram[55] = "m";
ram[56] = "?";
ram[57] = " ";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
18 : begin
ram[0] = "A";
ram[1] = " ";
ram[2] = "g";
ram[3] = "r";
ram[4] = "e";
ram[5] = "a";
ram[6] = "t";
ram[7] = " ";
ram[8] = "p";
ram[9] = "e";
ram[10] = "a";
ram[11] = "c";
ram[12] = "e";
ram[13] = " ";
ram[14] = "f";
ram[15] = "a";
ram[16] = "l";
ram[17] = "l";
ram[18] = "s";
ram[19] = " ";
ram[20] = "o";
ram[21] = "v";
ram[22] = "e";
ram[23] = "r";
ram[24] = " ";
ram[25] = "t";
ram[26] = "h";
ram[27] = "e";
ram[28] = " ";
ram[29] = "k";
ram[30] = "i";
ram[31] = "n";
ram[32] = "g";
ram[33] = "d";
ram[34] = "o";
ram[35] = "m";
ram[36] = ".";
ram[37] = " ";
ram[38] = "A";
ram[39] = "b";
ram[40] = "o";
ram[41] = "l";
ram[42] = "i";
ram[43] = "s";
ram[44] = "h";
ram[45] = " ";
ram[46] = "c";
ram[47] = "o";
ram[48] = "n";
ram[49] = "s";
ram[50] = "c";
ram[51] = "r";
ram[52] = "i";
ram[53] = "p";
ram[54] = "t";
ram[55] = "i";
ram[56] = "o";
ram[57] = "n";
ram[58] = "?";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
19 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "n";
ram[5] = "e";
ram[6] = "i";
ram[7] = "g";
ram[8] = "h";
ram[9] = "b";
ram[10] = "o";
ram[11] = "u";
ram[12] = "r";
ram[13] = "i";
ram[14] = "n";
ram[15] = "g";
ram[16] = " ";
ram[17] = "k";
ram[18] = "i";
ram[19] = "n";
ram[20] = "g";
ram[21] = " ";
ram[22] = "i";
ram[23] = "s";
ram[24] = " ";
ram[25] = "v";
ram[26] = "i";
ram[27] = "s";
ram[28] = "i";
ram[29] = "t";
ram[30] = "i";
ram[31] = "n";
ram[32] = "g";
ram[33] = ".";
ram[34] = " ";
ram[35] = "O";
ram[36] = "r";
ram[37] = "g";
ram[38] = "a";
ram[39] = "n";
ram[40] = "i";
ram[41] = "z";
ram[42] = "e";
ram[43] = " ";
ram[44] = "a";
ram[45] = " ";
ram[46] = "g";
ram[47] = "r";
ram[48] = "a";
ram[49] = "n";
ram[50] = "d";
ram[51] = " ";
ram[52] = "f";
ram[53] = "e";
ram[54] = "a";
ram[55] = "s";
ram[56] = "t";
ram[57] = "?";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
20 : begin
ram[0] = "O";
ram[1] = "u";
ram[2] = "r";
ram[3] = " ";
ram[4] = "w";
ram[5] = "e";
ram[6] = "a";
ram[7] = "p";
ram[8] = "o";
ram[9] = "n";
ram[10] = "r";
ram[11] = "y";
ram[12] = " ";
ram[13] = "i";
ram[14] = "s";
ram[15] = " ";
ram[16] = "o";
ram[17] = "u";
ram[18] = "t";
ram[19] = "d";
ram[20] = "a";
ram[21] = "t";
ram[22] = "e";
ram[23] = "d";
ram[24] = ".";
ram[25] = " ";
ram[26] = "I";
ram[27] = "n";
ram[28] = "v";
ram[29] = "e";
ram[30] = "s";
ram[31] = "t";
ram[32] = " ";
ram[33] = "i";
ram[34] = "n";
ram[35] = " ";
ram[36] = "s";
ram[37] = "p";
ram[38] = "o";
ram[39] = "o";
ram[40] = "n";
ram[41] = "s";
ram[42] = " ";
ram[43] = "t";
ram[44] = "o";
ram[45] = " ";
ram[46] = "m";
ram[47] = "a";
ram[48] = "k";
ram[49] = "e";
ram[50] = " ";
ram[51] = "o";
ram[52] = "u";
ram[53] = "r";
ram[54] = " ";
ram[55] = "w";
ram[56] = "e";
ram[57] = "a";
ram[58] = "p";
ram[59] = "o";
ram[60] = "n";
ram[61] = "s";
ram[62] = " ";
ram[63] = "s";
ram[64] = "t";
ram[65] = "r";
ram[66] = "o";
ram[67] = "n";
ram[68] = "g";
ram[69] = "e";
ram[70] = "r";
ram[71] = "?";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
21 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = "r";
ram[4] = "e";
ram[5] = " ";
ram[6] = "h";
ram[7] = "a";
ram[8] = "s";
ram[9] = " ";
ram[10] = "n";
ram[11] = "o";
ram[12] = "t";
ram[13] = " ";
ram[14] = "b";
ram[15] = "e";
ram[16] = "e";
ram[17] = "n";
ram[18] = " ";
ram[19] = "a";
ram[20] = " ";
ram[21] = "w";
ram[22] = "a";
ram[23] = "r";
ram[24] = " ";
ram[25] = "i";
ram[26] = "n";
ram[27] = " ";
ram[28] = "a";
ram[29] = "g";
ram[30] = "e";
ram[31] = "s";
ram[32] = ".";
ram[33] = " ";
ram[34] = "G";
ram[35] = "i";
ram[36] = "v";
ram[37] = "e";
ram[38] = " ";
ram[39] = "a";
ram[40] = " ";
ram[41] = "r";
ram[42] = "a";
ram[43] = "l";
ram[44] = "l";
ram[45] = "y";
ram[46] = "i";
ram[47] = "n";
ram[48] = "g";
ram[49] = " ";
ram[50] = "s";
ram[51] = "p";
ram[52] = "e";
ram[53] = "e";
ram[54] = "c";
ram[55] = "h";
ram[56] = " ";
ram[57] = "t";
ram[58] = "o";
ram[59] = " ";
ram[60] = "t";
ram[61] = "h";
ram[62] = "e";
ram[63] = " ";
ram[64] = "m";
ram[65] = "i";
ram[66] = "l";
ram[67] = "i";
ram[68] = "t";
ram[69] = "a";
ram[70] = "r";
ram[71] = "y";
ram[72] = "?";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
22 : begin
ram[0] = "Y";
ram[1] = "o";
ram[2] = "u";
ram[3] = "r";
ram[4] = " ";
ram[5] = "f";
ram[6] = "o";
ram[7] = "r";
ram[8] = "t";
ram[9] = "r";
ram[10] = "e";
ram[11] = "s";
ram[12] = "s";
ram[13] = " ";
ram[14] = "i";
ram[15] = "s";
ram[16] = " ";
ram[17] = "w";
ram[18] = "e";
ram[19] = "a";
ram[20] = "k";
ram[21] = ".";
ram[22] = " ";
ram[23] = "B";
ram[24] = "u";
ram[25] = "i";
ram[26] = "l";
ram[27] = "d";
ram[28] = " ";
ram[29] = "a";
ram[30] = "n";
ram[31] = "o";
ram[32] = "t";
ram[33] = "h";
ram[34] = "e";
ram[35] = "r";
ram[36] = " ";
ram[37] = "t";
ram[38] = "o";
ram[39] = "w";
ram[40] = "e";
ram[41] = "r";
ram[42] = "?";
ram[43] = " ";
ram[44] = " ";
ram[45] = " ";
ram[46] = " ";
ram[47] = " ";
ram[48] = " ";
ram[49] = " ";
ram[50] = " ";
ram[51] = " ";
ram[52] = " ";
ram[53] = " ";
ram[54] = " ";
ram[55] = " ";
ram[56] = " ";
ram[57] = " ";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
23 : begin
ram[0] = "Y";
ram[1] = "o";
ram[2] = "u";
ram[3] = "r";
ram[4] = " ";
ram[5] = "a";
ram[6] = "l";
ram[7] = "l";
ram[8] = "i";
ram[9] = "e";
ram[10] = "d";
ram[11] = " ";
ram[12] = "n";
ram[13] = "a";
ram[14] = "t";
ram[15] = "i";
ram[16] = "o";
ram[17] = "n";
ram[18] = "s";
ram[19] = " ";
ram[20] = "r";
ram[21] = "e";
ram[22] = "q";
ram[23] = "u";
ram[24] = "i";
ram[25] = "r";
ram[26] = "e";
ram[27] = " ";
ram[28] = "y";
ram[29] = "o";
ram[30] = "u";
ram[31] = "r";
ram[32] = " ";
ram[33] = "m";
ram[34] = "i";
ram[35] = "l";
ram[36] = "i";
ram[37] = "t";
ram[38] = "a";
ram[39] = "r";
ram[40] = "y";
ram[41] = " ";
ram[42] = "s";
ram[43] = "u";
ram[44] = "p";
ram[45] = "p";
ram[46] = "o";
ram[47] = "r";
ram[48] = "t";
ram[49] = ".";
ram[50] = " ";
ram[51] = "A";
ram[52] = "s";
ram[53] = "s";
ram[54] = "i";
ram[55] = "s";
ram[56] = "t";
ram[57] = " ";
ram[58] = "t";
ram[59] = "h";
ram[60] = "e";
ram[61] = "m";
ram[62] = "?";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
24 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = "r";
ram[4] = "e";
ram[5] = " ";
ram[6] = "h";
ram[7] = "a";
ram[8] = "s";
ram[9] = " ";
ram[10] = "b";
ram[11] = "e";
ram[12] = "e";
ram[13] = "n";
ram[14] = " ";
ram[15] = "a";
ram[16] = " ";
ram[17] = "b";
ram[18] = "a";
ram[19] = "d";
ram[20] = " ";
ram[21] = "h";
ram[22] = "a";
ram[23] = "r";
ram[24] = "v";
ram[25] = "e";
ram[26] = "s";
ram[27] = "t";
ram[28] = " ";
ram[29] = "t";
ram[30] = "h";
ram[31] = "i";
ram[32] = "s";
ram[33] = " ";
ram[34] = "s";
ram[35] = "e";
ram[36] = "a";
ram[37] = "s";
ram[38] = "o";
ram[39] = "n";
ram[40] = ".";
ram[41] = " ";
ram[42] = "D";
ram[43] = "e";
ram[44] = "c";
ram[45] = "r";
ram[46] = "e";
ram[47] = "a";
ram[48] = "s";
ram[49] = "e";
ram[50] = " ";
ram[51] = "t";
ram[52] = "a";
ram[53] = "x";
ram[54] = "e";
ram[55] = "s";
ram[56] = "?";
ram[57] = " ";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
25 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "p";
ram[5] = "e";
ram[6] = "o";
ram[7] = "p";
ram[8] = "l";
ram[9] = "e";
ram[10] = " ";
ram[11] = "f";
ram[12] = "e";
ram[13] = "e";
ram[14] = "l";
ram[15] = " ";
ram[16] = "t";
ram[17] = "h";
ram[18] = "a";
ram[19] = "t";
ram[20] = " ";
ram[21] = "t";
ram[22] = "h";
ram[23] = "e";
ram[24] = " ";
ram[25] = "p";
ram[26] = "r";
ram[27] = "i";
ram[28] = "c";
ram[29] = "e";
ram[30] = " ";
ram[31] = "o";
ram[32] = "f";
ram[33] = " ";
ram[34] = "b";
ram[35] = "r";
ram[36] = "e";
ram[37] = "a";
ram[38] = "d";
ram[39] = " ";
ram[40] = "i";
ram[41] = "s";
ram[42] = " ";
ram[43] = "t";
ram[44] = "o";
ram[45] = "o";
ram[46] = " ";
ram[47] = "h";
ram[48] = "i";
ram[49] = "g";
ram[50] = "h";
ram[51] = ".";
ram[52] = " ";
ram[53] = "L";
ram[54] = "o";
ram[55] = "w";
ram[56] = "e";
ram[57] = "r";
ram[58] = " ";
ram[59] = "t";
ram[60] = "h";
ram[61] = "e";
ram[62] = " ";
ram[63] = "p";
ram[64] = "r";
ram[65] = "i";
ram[66] = "c";
ram[67] = "e";
ram[68] = "?";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
26 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "s";
ram[5] = "t";
ram[6] = "r";
ram[7] = "e";
ram[8] = "e";
ram[9] = "t";
ram[10] = "s";
ram[11] = " ";
ram[12] = "s";
ram[13] = "m";
ram[14] = "e";
ram[15] = "l";
ram[16] = "l";
ram[17] = " ";
ram[18] = "l";
ram[19] = "i";
ram[20] = "k";
ram[21] = "e";
ram[22] = " ";
ram[23] = "s";
ram[24] = "e";
ram[25] = "w";
ram[26] = "a";
ram[27] = "g";
ram[28] = "e";
ram[29] = ".";
ram[30] = " ";
ram[31] = "C";
ram[32] = "l";
ram[33] = "e";
ram[34] = "a";
ram[35] = "r";
ram[36] = " ";
ram[37] = "t";
ram[38] = "h";
ram[39] = "e";
ram[40] = " ";
ram[41] = "s";
ram[42] = "e";
ram[43] = "w";
ram[44] = "a";
ram[45] = "g";
ram[46] = "e";
ram[47] = " ";
ram[48] = "s";
ram[49] = "y";
ram[50] = "s";
ram[51] = "t";
ram[52] = "e";
ram[53] = "m";
ram[54] = "?";
ram[55] = " ";
ram[56] = " ";
ram[57] = " ";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
27 : begin
ram[0] = "I";
ram[1] = "t";
ram[2] = " ";
ram[3] = "i";
ram[4] = "s";
ram[5] = " ";
ram[6] = "y";
ram[7] = "o";
ram[8] = "u";
ram[9] = "r";
ram[10] = " ";
ram[11] = "k";
ram[12] = "i";
ram[13] = "n";
ram[14] = "g";
ram[15] = "d";
ram[16] = "o";
ram[17] = "m";
ram[18] = "s";
ram[19] = " ";
ram[20] = "a";
ram[21] = "n";
ram[22] = "n";
ram[23] = "i";
ram[24] = "v";
ram[25] = "e";
ram[26] = "r";
ram[27] = "s";
ram[28] = "a";
ram[29] = "r";
ram[30] = "y";
ram[31] = ".";
ram[32] = " ";
ram[33] = "H";
ram[34] = "o";
ram[35] = "l";
ram[36] = "d";
ram[37] = " ";
ram[38] = "a";
ram[39] = " ";
ram[40] = "f";
ram[41] = "e";
ram[42] = "a";
ram[43] = "s";
ram[44] = "t";
ram[45] = " ";
ram[46] = "t";
ram[47] = "o";
ram[48] = " ";
ram[49] = "c";
ram[50] = "e";
ram[51] = "l";
ram[52] = "e";
ram[53] = "b";
ram[54] = "r";
ram[55] = "a";
ram[56] = "t";
ram[57] = "e";
ram[58] = "?";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
28 : begin
ram[0] = "Y";
ram[1] = "o";
ram[2] = "u";
ram[3] = "r";
ram[4] = " ";
ram[5] = "k";
ram[6] = "i";
ram[7] = "n";
ram[8] = "g";
ram[9] = "d";
ram[10] = "o";
ram[11] = "m";
ram[12] = " ";
ram[13] = "f";
ram[14] = "i";
ram[15] = "n";
ram[16] = "a";
ram[17] = "n";
ram[18] = "c";
ram[19] = "e";
ram[20] = "s";
ram[21] = " ";
ram[22] = "a";
ram[23] = "r";
ram[24] = "e";
ram[25] = " ";
ram[26] = "l";
ram[27] = "o";
ram[28] = "w";
ram[29] = ".";
ram[30] = " ";
ram[31] = "S";
ram[32] = "t";
ram[33] = "a";
ram[34] = "r";
ram[35] = "t";
ram[36] = " ";
ram[37] = "a";
ram[38] = " ";
ram[39] = "p";
ram[40] = "y";
ram[41] = "r";
ram[42] = "a";
ram[43] = "m";
ram[44] = "i";
ram[45] = "d";
ram[46] = " ";
ram[47] = "s";
ram[48] = "c";
ram[49] = "h";
ram[50] = "e";
ram[51] = "m";
ram[52] = "e";
ram[53] = "?";
ram[54] = " ";
ram[55] = " ";
ram[56] = " ";
ram[57] = " ";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
29 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "p";
ram[5] = "r";
ram[6] = "i";
ram[7] = "e";
ram[8] = "s";
ram[9] = "t";
ram[10] = "s";
ram[11] = " ";
ram[12] = "w";
ram[13] = "o";
ram[14] = "u";
ram[15] = "l";
ram[16] = "d";
ram[17] = " ";
ram[18] = "l";
ram[19] = "i";
ram[20] = "k";
ram[21] = "e";
ram[22] = " ";
ram[23] = "t";
ram[24] = "o";
ram[25] = " ";
ram[26] = "h";
ram[27] = "o";
ram[28] = "l";
ram[29] = "d";
ram[30] = " ";
ram[31] = "a";
ram[32] = " ";
ram[33] = "m";
ram[34] = "a";
ram[35] = "s";
ram[36] = "s";
ram[37] = " ";
ram[38] = "p";
ram[39] = "r";
ram[40] = "a";
ram[41] = "y";
ram[42] = "e";
ram[43] = "r";
ram[44] = ".";
ram[45] = " ";
ram[46] = "A";
ram[47] = "l";
ram[48] = "l";
ram[49] = "o";
ram[50] = "w";
ram[51] = " ";
ram[52] = "t";
ram[53] = "h";
ram[54] = "e";
ram[55] = "m";
ram[56] = " ";
ram[57] = "t";
ram[58] = "o";
ram[59] = " ";
ram[60] = "p";
ram[61] = "r";
ram[62] = "o";
ram[63] = "c";
ram[64] = "e";
ram[65] = "e";
ram[66] = "d";
ram[67] = "?";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
30 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "p";
ram[5] = "r";
ram[6] = "i";
ram[7] = "e";
ram[8] = "s";
ram[9] = "t";
ram[10] = " ";
ram[11] = "d";
ram[12] = "e";
ram[13] = "f";
ram[14] = "e";
ram[15] = "c";
ram[16] = "a";
ram[17] = "t";
ram[18] = "e";
ram[19] = "d";
ram[20] = " ";
ram[21] = "o";
ram[22] = "n";
ram[23] = " ";
ram[24] = "y";
ram[25] = "o";
ram[26] = "u";
ram[27] = "r";
ram[28] = " ";
ram[29] = "d";
ram[30] = "o";
ram[31] = "o";
ram[32] = "r";
ram[33] = "s";
ram[34] = "t";
ram[35] = "e";
ram[36] = "p";
ram[37] = ".";
ram[38] = " ";
ram[39] = "S";
ram[40] = "t";
ram[41] = "a";
ram[42] = "r";
ram[43] = "t";
ram[44] = " ";
ram[45] = "a";
ram[46] = " ";
ram[47] = "c";
ram[48] = "u";
ram[49] = "l";
ram[50] = "t";
ram[51] = "?";
ram[52] = " ";
ram[53] = " ";
ram[54] = " ";
ram[55] = " ";
ram[56] = " ";
ram[57] = " ";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
31 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "g";
ram[5] = "e";
ram[6] = "n";
ram[7] = "e";
ram[8] = "r";
ram[9] = "a";
ram[10] = "l";
ram[11] = " ";
ram[12] = "w";
ram[13] = "a";
ram[14] = "n";
ram[15] = "t";
ram[16] = "s";
ram[17] = " ";
ram[18] = "t";
ram[19] = "o";
ram[20] = " ";
ram[21] = "d";
ram[22] = "e";
ram[23] = "m";
ram[24] = "o";
ram[25] = "n";
ram[26] = "s";
ram[27] = "t";
ram[28] = "r";
ram[29] = "a";
ram[30] = "t";
ram[31] = "e";
ram[32] = " ";
ram[33] = "h";
ram[34] = "i";
ram[35] = "s";
ram[36] = " ";
ram[37] = "m";
ram[38] = "e";
ram[39] = "n";
ram[40] = "'";
ram[41] = "s";
ram[42] = " ";
ram[43] = "p";
ram[44] = "r";
ram[45] = "o";
ram[46] = "w";
ram[47] = "e";
ram[48] = "s";
ram[49] = "s";
ram[50] = ".";
ram[51] = " ";
ram[52] = "A";
ram[53] = "c";
ram[54] = "c";
ram[55] = "e";
ram[56] = "p";
ram[57] = "t";
ram[58] = "?";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
32 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "g";
ram[5] = "e";
ram[6] = "n";
ram[7] = "e";
ram[8] = "r";
ram[9] = "a";
ram[10] = "l";
ram[11] = " ";
ram[12] = "w";
ram[13] = "a";
ram[14] = "n";
ram[15] = "t";
ram[16] = "s";
ram[17] = " ";
ram[18] = "t";
ram[19] = "o";
ram[20] = " ";
ram[21] = "y";
ram[22] = "o";
ram[23] = "u";
ram[24] = " ";
ram[25] = "t";
ram[26] = "o";
ram[27] = " ";
ram[28] = "i";
ram[29] = "n";
ram[30] = "s";
ram[31] = "p";
ram[32] = "e";
ram[33] = "c";
ram[34] = "t";
ram[35] = " ";
ram[36] = "h";
ram[37] = "i";
ram[38] = "s";
ram[39] = " ";
ram[40] = "c";
ram[41] = "a";
ram[42] = "n";
ram[43] = "n";
ram[44] = "o";
ram[45] = "n";
ram[46] = "s";
ram[47] = ".";
ram[48] = " ";
ram[49] = "W";
ram[50] = "e";
ram[51] = "a";
ram[52] = "r";
ram[53] = " ";
ram[54] = "g";
ram[55] = "l";
ram[56] = "o";
ram[57] = "v";
ram[58] = "e";
ram[59] = "s";
ram[60] = "?";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
33 : begin
ram[0] = "B";
ram[1] = "e";
ram[2] = "g";
ram[3] = "g";
ram[4] = "a";
ram[5] = "r";
ram[6] = "s";
ram[7] = " ";
ram[8] = "a";
ram[9] = "r";
ram[10] = "e";
ram[11] = " ";
ram[12] = "i";
ram[13] = "n";
ram[14] = "v";
ram[15] = "a";
ram[16] = "d";
ram[17] = "i";
ram[18] = "n";
ram[19] = "g";
ram[20] = " ";
ram[21] = "t";
ram[22] = "h";
ram[23] = "e";
ram[24] = " ";
ram[25] = "s";
ram[26] = "t";
ram[27] = "r";
ram[28] = "e";
ram[29] = "e";
ram[30] = "t";
ram[31] = "s";
ram[32] = ".";
ram[33] = " ";
ram[34] = "T";
ram[35] = "h";
ram[36] = "r";
ram[37] = "o";
ram[38] = "w";
ram[39] = " ";
ram[40] = "t";
ram[41] = "h";
ram[42] = "e";
ram[43] = "m";
ram[44] = " ";
ram[45] = "o";
ram[46] = "u";
ram[47] = "t";
ram[48] = "?";
ram[49] = " ";
ram[50] = " ";
ram[51] = " ";
ram[52] = " ";
ram[53] = " ";
ram[54] = " ";
ram[55] = " ";
ram[56] = " ";
ram[57] = " ";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
34 : begin
ram[0] = "A";
ram[1] = " ";
ram[2] = "h";
ram[3] = "u";
ram[4] = "n";
ram[5] = "g";
ram[6] = "r";
ram[7] = "y";
ram[8] = " ";
ram[9] = "b";
ram[10] = "o";
ram[11] = "y";
ram[12] = " ";
ram[13] = "w";
ram[14] = "a";
ram[15] = "s";
ram[16] = " ";
ram[17] = "c";
ram[18] = "a";
ram[19] = "u";
ram[20] = "g";
ram[21] = "h";
ram[22] = "t";
ram[23] = " ";
ram[24] = "s";
ram[25] = "t";
ram[26] = "e";
ram[27] = "a";
ram[28] = "l";
ram[29] = "i";
ram[30] = "n";
ram[31] = "g";
ram[32] = " ";
ram[33] = "y";
ram[34] = "o";
ram[35] = "u";
ram[36] = "r";
ram[37] = " ";
ram[38] = "c";
ram[39] = "r";
ram[40] = "o";
ram[41] = "w";
ram[42] = "n";
ram[43] = " ";
ram[44] = "j";
ram[45] = "e";
ram[46] = "w";
ram[47] = "e";
ram[48] = "l";
ram[49] = "s";
ram[50] = ".";
ram[51] = " ";
ram[52] = "B";
ram[53] = "r";
ram[54] = "i";
ram[55] = "n";
ram[56] = "g";
ram[57] = " ";
ram[58] = "h";
ram[59] = "i";
ram[60] = "m";
ram[61] = " ";
ram[62] = "t";
ram[63] = "o";
ram[64] = " ";
ram[65] = "t";
ram[66] = "h";
ram[67] = "e";
ram[68] = " ";
ram[69] = "p";
ram[70] = "r";
ram[71] = "i";
ram[72] = "e";
ram[73] = "s";
ram[74] = "t";
ram[75] = "?";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
35 : begin
ram[0] = "K";
ram[1] = "i";
ram[2] = "n";
ram[3] = "g";
ram[4] = "d";
ram[5] = "o";
ram[6] = "m";
ram[7] = "s";
ram[8] = " ";
ram[9] = "f";
ram[10] = "r";
ram[11] = "o";
ram[12] = "m";
ram[13] = " ";
ram[14] = "t";
ram[15] = "h";
ram[16] = "e";
ram[17] = " ";
ram[18] = "o";
ram[19] = "r";
ram[20] = "i";
ram[21] = "e";
ram[22] = "n";
ram[23] = "t";
ram[24] = " ";
ram[25] = "w";
ram[26] = "o";
ram[27] = "u";
ram[28] = "l";
ram[29] = "d";
ram[30] = " ";
ram[31] = "l";
ram[32] = "i";
ram[33] = "k";
ram[34] = "e";
ram[35] = " ";
ram[36] = "t";
ram[37] = "o";
ram[38] = " ";
ram[39] = "s";
ram[40] = "i";
ram[41] = "g";
ram[42] = "n";
ram[43] = " ";
ram[44] = "a";
ram[45] = " ";
ram[46] = "t";
ram[47] = "r";
ram[48] = "a";
ram[49] = "d";
ram[50] = "e";
ram[51] = " ";
ram[52] = "p";
ram[53] = "a";
ram[54] = "c";
ram[55] = "t";
ram[56] = ".";
ram[57] = " ";
ram[58] = "S";
ram[59] = "i";
ram[60] = "g";
ram[61] = "n";
ram[62] = " ";
ram[63] = "t";
ram[64] = "h";
ram[65] = "e";
ram[66] = " ";
ram[67] = "t";
ram[68] = "r";
ram[69] = "e";
ram[70] = "a";
ram[71] = "t";
ram[72] = "y";
ram[73] = "?";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
36 : begin
ram[0] = "Y";
ram[1] = "o";
ram[2] = "u";
ram[3] = "r";
ram[4] = " ";
ram[5] = "n";
ram[6] = "o";
ram[7] = "r";
ram[8] = "t";
ram[9] = "h";
ram[10] = "e";
ram[11] = "r";
ram[12] = "n";
ram[13] = " ";
ram[14] = "n";
ram[15] = "e";
ram[16] = "i";
ram[17] = "g";
ram[18] = "h";
ram[19] = "b";
ram[20] = "o";
ram[21] = "u";
ram[22] = "r";
ram[23] = "s";
ram[24] = " ";
ram[25] = "w";
ram[26] = "a";
ram[27] = "n";
ram[28] = "t";
ram[29] = " ";
ram[30] = "y";
ram[31] = "o";
ram[32] = "u";
ram[33] = " ";
ram[34] = "t";
ram[35] = "o";
ram[36] = " ";
ram[37] = "p";
ram[38] = "a";
ram[39] = "y";
ram[40] = " ";
ram[41] = "f";
ram[42] = "o";
ram[43] = "r";
ram[44] = " ";
ram[45] = "t";
ram[46] = "h";
ram[47] = "e";
ram[48] = "i";
ram[49] = "r";
ram[50] = " ";
ram[51] = "b";
ram[52] = "o";
ram[53] = "r";
ram[54] = "d";
ram[55] = "e";
ram[56] = "r";
ram[57] = " ";
ram[58] = "w";
ram[59] = "a";
ram[60] = "l";
ram[61] = "l";
ram[62] = ".";
ram[63] = " ";
ram[64] = "S";
ram[65] = "i";
ram[66] = "?";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
37 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "h";
ram[5] = "e";
ram[6] = "a";
ram[7] = "d";
ram[8] = " ";
ram[9] = "p";
ram[10] = "r";
ram[11] = "i";
ram[12] = "e";
ram[13] = "s";
ram[14] = "t";
ram[15] = " ";
ram[16] = "h";
ram[17] = "a";
ram[18] = "s";
ram[19] = " ";
ram[20] = "b";
ram[21] = "e";
ram[22] = "c";
ram[23] = "o";
ram[24] = "m";
ram[25] = "e";
ram[26] = " ";
ram[27] = "t";
ram[28] = "o";
ram[29] = "o";
ram[30] = " ";
ram[31] = "o";
ram[32] = "l";
ram[33] = "d";
ram[34] = " ";
ram[35] = "a";
ram[36] = "n";
ram[37] = "d";
ram[38] = " ";
ram[39] = "h";
ram[40] = "a";
ram[41] = "s";
ram[42] = " ";
ram[43] = "r";
ram[44] = "e";
ram[45] = "t";
ram[46] = "i";
ram[47] = "r";
ram[48] = "e";
ram[49] = "d";
ram[50] = ",";
ram[51] = " ";
ram[52] = "t";
ram[53] = "h";
ram[54] = "e";
ram[55] = " ";
ram[56] = "c";
ram[57] = "h";
ram[58] = "u";
ram[59] = "r";
ram[60] = "c";
ram[61] = "h";
ram[62] = " ";
ram[63] = "i";
ram[64] = "s";
ram[65] = " ";
ram[66] = "u";
ram[67] = "n";
ram[68] = "s";
ram[69] = "t";
ram[70] = "a";
ram[71] = "b";
ram[72] = "l";
ram[73] = "e";
ram[74] = ".";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
38 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "p";
ram[5] = "e";
ram[6] = "o";
ram[7] = "p";
ram[8] = "l";
ram[9] = "e";
ram[10] = " ";
ram[11] = "a";
ram[12] = "r";
ram[13] = "e";
ram[14] = " ";
ram[15] = "h";
ram[16] = "a";
ram[17] = "p";
ram[18] = "p";
ram[19] = "y";
ram[20] = " ";
ram[21] = "a";
ram[22] = "n";
ram[23] = "d";
ram[24] = " ";
ram[25] = "y";
ram[26] = "o";
ram[27] = "u";
ram[28] = " ";
ram[29] = "a";
ram[30] = "r";
ram[31] = "e";
ram[32] = " ";
ram[33] = "l";
ram[34] = "o";
ram[35] = "v";
ram[36] = "e";
ram[37] = "d";
ram[38] = " ";
ram[39] = "b";
ram[40] = "y";
ram[41] = " ";
ram[42] = "t";
ram[43] = "h";
ram[44] = "e";
ram[45] = "m";
ram[46] = ".";
ram[47] = " ";
ram[48] = " ";
ram[49] = " ";
ram[50] = " ";
ram[51] = " ";
ram[52] = " ";
ram[53] = " ";
ram[54] = " ";
ram[55] = " ";
ram[56] = " ";
ram[57] = " ";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
39 : begin
ram[0] = "A";
ram[1] = " ";
ram[2] = "m";
ram[3] = "e";
ram[4] = "t";
ram[5] = "e";
ram[6] = "o";
ram[7] = "r";
ram[8] = " ";
ram[9] = "d";
ram[10] = "e";
ram[11] = "s";
ram[12] = "t";
ram[13] = "r";
ram[14] = "o";
ram[15] = "y";
ram[16] = "e";
ram[17] = "d";
ram[18] = " ";
ram[19] = "t";
ram[20] = "h";
ram[21] = "e";
ram[22] = " ";
ram[23] = "n";
ram[24] = "e";
ram[25] = "i";
ram[26] = "g";
ram[27] = "h";
ram[28] = "b";
ram[29] = "o";
ram[30] = "u";
ram[31] = "r";
ram[32] = "i";
ram[33] = "n";
ram[34] = "g";
ram[35] = " ";
ram[36] = "c";
ram[37] = "i";
ram[38] = "t";
ram[39] = "y";
ram[40] = "!";
ram[41] = " ";
ram[42] = " ";
ram[43] = " ";
ram[44] = " ";
ram[45] = " ";
ram[46] = " ";
ram[47] = " ";
ram[48] = " ";
ram[49] = " ";
ram[50] = " ";
ram[51] = " ";
ram[52] = " ";
ram[53] = " ";
ram[54] = " ";
ram[55] = " ";
ram[56] = " ";
ram[57] = " ";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
40 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "p";
ram[5] = "r";
ram[6] = "e";
ram[7] = "v";
ram[8] = "i";
ram[9] = "o";
ram[10] = "u";
ram[11] = "s";
ram[12] = " ";
ram[13] = "K";
ram[14] = "i";
ram[15] = "n";
ram[16] = "g";
ram[17] = " ";
ram[18] = "t";
ram[19] = "o";
ram[20] = "o";
ram[21] = "k";
ram[22] = " ";
ram[23] = "a";
ram[24] = " ";
ram[25] = "l";
ram[26] = "o";
ram[27] = "a";
ram[28] = "n";
ram[29] = " ";
ram[30] = "a";
ram[31] = "n";
ram[32] = "d";
ram[33] = " ";
ram[34] = "n";
ram[35] = "o";
ram[36] = "w";
ram[37] = " ";
ram[38] = "t";
ram[39] = "h";
ram[40] = "e";
ram[41] = " ";
ram[42] = "d";
ram[43] = "e";
ram[44] = "b";
ram[45] = "t";
ram[46] = " ";
ram[47] = "m";
ram[48] = "u";
ram[49] = "s";
ram[50] = "t";
ram[51] = " ";
ram[52] = "b";
ram[53] = "e";
ram[54] = " ";
ram[55] = "r";
ram[56] = "e";
ram[57] = "p";
ram[58] = "a";
ram[59] = "i";
ram[60] = "d";
ram[61] = ".";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
41 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "k";
ram[5] = "i";
ram[6] = "n";
ram[7] = "g";
ram[8] = "d";
ram[9] = "o";
ram[10] = "m";
ram[11] = "s";
ram[12] = " ";
ram[13] = "i";
ram[14] = "n";
ram[15] = " ";
ram[16] = "t";
ram[17] = "h";
ram[18] = "e";
ram[19] = " ";
ram[20] = "o";
ram[21] = "r";
ram[22] = "i";
ram[23] = "e";
ram[24] = "n";
ram[25] = "t";
ram[26] = " ";
ram[27] = "h";
ram[28] = "a";
ram[29] = "v";
ram[30] = "e";
ram[31] = " ";
ram[32] = "s";
ram[33] = "e";
ram[34] = "i";
ram[35] = "z";
ram[36] = "e";
ram[37] = "d";
ram[38] = " ";
ram[39] = "y";
ram[40] = "o";
ram[41] = "u";
ram[42] = "r";
ram[43] = " ";
ram[44] = "t";
ram[45] = "r";
ram[46] = "e";
ram[47] = "b";
ram[48] = "u";
ram[49] = "c";
ram[50] = "h";
ram[51] = "e";
ram[52] = "t";
ram[53] = "s";
ram[54] = ".";
ram[55] = " ";
ram[56] = " ";
ram[57] = " ";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
42 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "n";
ram[5] = "e";
ram[6] = "i";
ram[7] = "g";
ram[8] = "h";
ram[9] = "b";
ram[10] = "o";
ram[11] = "u";
ram[12] = "r";
ram[13] = "i";
ram[14] = "n";
ram[15] = "g";
ram[16] = " ";
ram[17] = "p";
ram[18] = "r";
ram[19] = "i";
ram[20] = "n";
ram[21] = "c";
ram[22] = "e";
ram[23] = " ";
ram[24] = "w";
ram[25] = "a";
ram[26] = "n";
ram[27] = "t";
ram[28] = "s";
ram[29] = " ";
ram[30] = "t";
ram[31] = "o";
ram[32] = " ";
ram[33] = "m";
ram[34] = "a";
ram[35] = "r";
ram[36] = "r";
ram[37] = "y";
ram[38] = " ";
ram[39] = "y";
ram[40] = "o";
ram[41] = "u";
ram[42] = "r";
ram[43] = " ";
ram[44] = "d";
ram[45] = "a";
ram[46] = "u";
ram[47] = "g";
ram[48] = "h";
ram[49] = "t";
ram[50] = "e";
ram[51] = "r";
ram[52] = ".";
ram[53] = " ";
ram[54] = "M";
ram[55] = "a";
ram[56] = "r";
ram[57] = "r";
ram[58] = "y";
ram[59] = " ";
ram[60] = "h";
ram[61] = "e";
ram[62] = "r";
ram[63] = " ";
ram[64] = "o";
ram[65] = "f";
ram[66] = "f";
ram[67] = "?";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
43 : begin
ram[0] = "R";
ram[1] = "e";
ram[2] = "l";
ram[3] = "a";
ram[4] = "t";
ram[5] = "i";
ram[6] = "o";
ram[7] = "n";
ram[8] = "s";
ram[9] = " ";
ram[10] = "w";
ram[11] = "i";
ram[12] = "t";
ram[13] = "h";
ram[14] = " ";
ram[15] = "t";
ram[16] = "h";
ram[17] = "e";
ram[18] = " ";
ram[19] = "n";
ram[20] = "e";
ram[21] = "i";
ram[22] = "g";
ram[23] = "h";
ram[24] = "b";
ram[25] = "o";
ram[26] = "u";
ram[27] = "r";
ram[28] = "i";
ram[29] = "n";
ram[30] = "g";
ram[31] = " ";
ram[32] = "k";
ram[33] = "i";
ram[34] = "n";
ram[35] = "g";
ram[36] = "d";
ram[37] = "o";
ram[38] = "m";
ram[39] = " ";
ram[40] = "a";
ram[41] = "r";
ram[42] = "e";
ram[43] = " ";
ram[44] = "d";
ram[45] = "e";
ram[46] = "t";
ram[47] = "e";
ram[48] = "r";
ram[49] = "i";
ram[50] = "o";
ram[51] = "r";
ram[52] = "a";
ram[53] = "t";
ram[54] = "i";
ram[55] = "n";
ram[56] = "g";
ram[57] = ".";
ram[58] = " ";
ram[59] = "S";
ram[60] = "e";
ram[61] = "n";
ram[62] = "d";
ram[63] = " ";
ram[64] = "g";
ram[65] = "i";
ram[66] = "f";
ram[67] = "t";
ram[68] = "s";
ram[69] = "?";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
44 : begin
ram[0] = "A";
ram[1] = " ";
ram[2] = "c";
ram[3] = "r";
ram[4] = "o";
ram[5] = "w";
ram[6] = " ";
ram[7] = "h";
ram[8] = "a";
ram[9] = "s";
ram[10] = " ";
ram[11] = "b";
ram[12] = "e";
ram[13] = "e";
ram[14] = "n";
ram[15] = " ";
ram[16] = "s";
ram[17] = "i";
ram[18] = "t";
ram[19] = "t";
ram[20] = "i";
ram[21] = "n";
ram[22] = "g";
ram[23] = " ";
ram[24] = "o";
ram[25] = "n";
ram[26] = " ";
ram[27] = "y";
ram[28] = "o";
ram[29] = "u";
ram[30] = "r";
ram[31] = " ";
ram[32] = "p";
ram[33] = "o";
ram[34] = "r";
ram[35] = "c";
ram[36] = "h";
ram[37] = " ";
ram[38] = "e";
ram[39] = "v";
ram[40] = "e";
ram[41] = "r";
ram[42] = "y";
ram[43] = " ";
ram[44] = "m";
ram[45] = "o";
ram[46] = "r";
ram[47] = "n";
ram[48] = "i";
ram[49] = "n";
ram[50] = "g";
ram[51] = ".";
ram[52] = " ";
ram[53] = "I";
ram[54] = "n";
ram[55] = "c";
ram[56] = "r";
ram[57] = "e";
ram[58] = "a";
ram[59] = "s";
ram[60] = "e";
ram[61] = " ";
ram[62] = "p";
ram[63] = "a";
ram[64] = "t";
ram[65] = "r";
ram[66] = "o";
ram[67] = "l";
ram[68] = "s";
ram[69] = "?";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
45 : begin
ram[0] = "Y";
ram[1] = "o";
ram[2] = "u";
ram[3] = " ";
ram[4] = "h";
ram[5] = "e";
ram[6] = "a";
ram[7] = "r";
ram[8] = " ";
ram[9] = "y";
ram[10] = "o";
ram[11] = "u";
ram[12] = "r";
ram[13] = " ";
ram[14] = "y";
ram[15] = "o";
ram[16] = "u";
ram[17] = "n";
ram[18] = "g";
ram[19] = "e";
ram[20] = "r";
ram[21] = " ";
ram[22] = "b";
ram[23] = "r";
ram[24] = "o";
ram[25] = "t";
ram[26] = "h";
ram[27] = "e";
ram[28] = "r";
ram[29] = " ";
ram[30] = "i";
ram[31] = "s";
ram[32] = " ";
ram[33] = "e";
ram[34] = "y";
ram[35] = "e";
ram[36] = "i";
ram[37] = "n";
ram[38] = "g";
ram[39] = " ";
ram[40] = "y";
ram[41] = "o";
ram[42] = "u";
ram[43] = "r";
ram[44] = " ";
ram[45] = "t";
ram[46] = "h";
ram[47] = "r";
ram[48] = "o";
ram[49] = "n";
ram[50] = "e";
ram[51] = ".";
ram[52] = " ";
ram[53] = "S";
ram[54] = "e";
ram[55] = "n";
ram[56] = "d";
ram[57] = " ";
ram[58] = "i";
ram[59] = "n";
ram[60] = "t";
ram[61] = "o";
ram[62] = " ";
ram[63] = "e";
ram[64] = "x";
ram[65] = "i";
ram[66] = "l";
ram[67] = "e";
ram[68] = "?";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
46 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "d";
ram[5] = "e";
ram[6] = "v";
ram[7] = "i";
ram[8] = "l";
ram[9] = " ";
ram[10] = "w";
ram[11] = "o";
ram[12] = "u";
ram[13] = "l";
ram[14] = "d";
ram[15] = " ";
ram[16] = "l";
ram[17] = "i";
ram[18] = "k";
ram[19] = "e";
ram[20] = " ";
ram[21] = "t";
ram[22] = "o";
ram[23] = " ";
ram[24] = "m";
ram[25] = "a";
ram[26] = "k";
ram[27] = "e";
ram[28] = " ";
ram[29] = "a";
ram[30] = " ";
ram[31] = "d";
ram[32] = "e";
ram[33] = "a";
ram[34] = "l";
ram[35] = " ";
ram[36] = "w";
ram[37] = "i";
ram[38] = "t";
ram[39] = "h";
ram[40] = " ";
ram[41] = "y";
ram[42] = "o";
ram[43] = "u";
ram[44] = ".";
ram[45] = " ";
ram[46] = " ";
ram[47] = " ";
ram[48] = " ";
ram[49] = " ";
ram[50] = " ";
ram[51] = " ";
ram[52] = " ";
ram[53] = " ";
ram[54] = " ";
ram[55] = " ";
ram[56] = " ";
ram[57] = " ";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
47 : begin
ram[0] = "D";
ram[1] = "i";
ram[2] = "j";
ram[3] = "k";
ram[4] = "s";
ram[5] = "t";
ram[6] = "r";
ram[7] = "a";
ram[8] = " ";
ram[9] = "t";
ram[10] = "h";
ram[11] = "e";
ram[12] = " ";
ram[13] = "S";
ram[14] = "h";
ram[15] = "o";
ram[16] = "r";
ram[17] = "t";
ram[18] = " ";
ram[19] = "w";
ram[20] = "a";
ram[21] = "s";
ram[22] = " ";
ram[23] = "c";
ram[24] = "a";
ram[25] = "u";
ram[26] = "g";
ram[27] = "h";
ram[28] = "t";
ram[29] = " ";
ram[30] = "t";
ram[31] = "r";
ram[32] = "e";
ram[33] = "s";
ram[34] = "p";
ram[35] = "a";
ram[36] = "s";
ram[37] = "s";
ram[38] = "i";
ram[39] = "n";
ram[40] = "g";
ram[41] = ".";
ram[42] = " ";
ram[43] = "Y";
ram[44] = "o";
ram[45] = "u";
ram[46] = "r";
ram[47] = " ";
ram[48] = "r";
ram[49] = "e";
ram[50] = "m";
ram[51] = "o";
ram[52] = "v";
ram[53] = "e";
ram[54] = " ";
ram[55] = "h";
ram[56] = "i";
ram[57] = "m";
ram[58] = " ";
ram[59] = "f";
ram[60] = "r";
ram[61] = "o";
ram[62] = "m";
ram[63] = " ";
ram[64] = "y";
ram[65] = "o";
ram[66] = "u";
ram[67] = "r";
ram[68] = " ";
ram[69] = "s";
ram[70] = "t";
ram[71] = "a";
ram[72] = "c";
ram[73] = "k";
ram[74] = ".";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
48 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "g";
ram[5] = "r";
ram[6] = "e";
ram[7] = "a";
ram[8] = "t";
ram[9] = " ";
ram[10] = "p";
ram[11] = "r";
ram[12] = "o";
ram[13] = "p";
ram[14] = "h";
ram[15] = "e";
ram[16] = "t";
ram[17] = " ";
ram[18] = "K";
ram[19] = "u";
ram[20] = "r";
ram[21] = "n";
ram[22] = "i";
ram[23] = "a";
ram[24] = "w";
ram[25] = "a";
ram[26] = "n";
ram[27] = " ";
ram[28] = "s";
ram[29] = "m";
ram[30] = "i";
ram[31] = "l";
ram[32] = "e";
ram[33] = "s";
ram[34] = " ";
ram[35] = "u";
ram[36] = "p";
ram[37] = "o";
ram[38] = "n";
ram[39] = " ";
ram[40] = "y";
ram[41] = "o";
ram[42] = "u";
ram[43] = ".";
ram[44] = " ";
ram[45] = " ";
ram[46] = " ";
ram[47] = " ";
ram[48] = " ";
ram[49] = " ";
ram[50] = " ";
ram[51] = " ";
ram[52] = " ";
ram[53] = " ";
ram[54] = " ";
ram[55] = " ";
ram[56] = " ";
ram[57] = " ";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
49 : begin
ram[0] = "A";
ram[1] = "d";
ram[2] = "v";
ram[3] = "i";
ram[4] = "s";
ram[5] = "o";
ram[6] = "r";
ram[7] = " ";
ram[8] = "Z";
ram[9] = "h";
ram[10] = "a";
ram[11] = "n";
ram[12] = "g";
ram[13] = " ";
ram[14] = "h";
ram[15] = "a";
ram[16] = "n";
ram[17] = "d";
ram[18] = "s";
ram[19] = " ";
ram[20] = "y";
ram[21] = "o";
ram[22] = "u";
ram[23] = " ";
ram[24] = "h";
ram[25] = "i";
ram[26] = "s";
ram[27] = " ";
ram[28] = "s";
ram[29] = "c";
ram[30] = "r";
ram[31] = "o";
ram[32] = "l";
ram[33] = "l";
ram[34] = "s";
ram[35] = " ";
ram[36] = "o";
ram[37] = "f";
ram[38] = " ";
ram[39] = "w";
ram[40] = "i";
ram[41] = "s";
ram[42] = "d";
ram[43] = "o";
ram[44] = "m";
ram[45] = ".";
ram[46] = " ";
ram[47] = " ";
ram[48] = " ";
ram[49] = " ";
ram[50] = " ";
ram[51] = " ";
ram[52] = " ";
ram[53] = " ";
ram[54] = " ";
ram[55] = " ";
ram[56] = " ";
ram[57] = " ";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
50 : begin
ram[0] = "I";
ram[1] = " ";
ram[2] = "A";
ram[3] = "M";
ram[4] = " ";
ram[5] = "A";
ram[6] = " ";
ram[7] = "F";
ram[8] = "I";
ram[9] = "L";
ram[10] = "E";
ram[11] = " ";
ram[12] = "A";
ram[13] = "N";
ram[14] = "D";
ram[15] = " ";
ram[16] = "Y";
ram[17] = "O";
ram[18] = "U";
ram[19] = " ";
ram[20] = "P";
ram[21] = "U";
ram[22] = "T";
ram[23] = " ";
ram[24] = "D";
ram[25] = "O";
ram[26] = "C";
ram[27] = "U";
ram[28] = "M";
ram[29] = "E";
ram[30] = "N";
ram[31] = "T";
ram[32] = "S";
ram[33] = " ";
ram[34] = "I";
ram[35] = "N";
ram[36] = " ";
ram[37] = "M";
ram[38] = "E";
ram[39] = ".";
ram[40] = "I";
ram[41] = " ";
ram[42] = "A";
ram[43] = "M";
ram[44] = " ";
ram[45] = "A";
ram[46] = " ";
ram[47] = "F";
ram[48] = "I";
ram[49] = "L";
ram[50] = "E";
ram[51] = " ";
ram[52] = "A";
ram[53] = "N";
ram[54] = "D";
ram[55] = " ";
ram[56] = "Y";
ram[57] = "O";
ram[58] = "U";
ram[59] = " ";
ram[60] = "P";
ram[61] = "U";
ram[62] = "T";
ram[63] = " ";
ram[64] = "D";
ram[65] = "O";
ram[66] = "C";
ram[67] = "U";
ram[68] = "M";
ram[69] = "E";
ram[70] = "N";
ram[71] = "T";
ram[72] = "S";
ram[73] = " ";
ram[74] = "I";
ram[75] = "N";
ram[76] = " ";
ram[77] = "M";
ram[78] = "E";
ram[79] = ".";
end
51 : begin
ram[0] = "Y";
ram[1] = "o";
ram[2] = "u";
ram[3] = "r";
ram[4] = " ";
ram[5] = "l";
ram[6] = "a";
ram[7] = "v";
ram[8] = "i";
ram[9] = "s";
ram[10] = "h";
ram[11] = " ";
ram[12] = "p";
ram[13] = "a";
ram[14] = "r";
ram[15] = "t";
ram[16] = "i";
ram[17] = "e";
ram[18] = "s";
ram[19] = " ";
ram[20] = "l";
ram[21] = "e";
ram[22] = "a";
ram[23] = "v";
ram[24] = "e";
ram[25] = " ";
ram[26] = "y";
ram[27] = "o";
ram[28] = "u";
ram[29] = " ";
ram[30] = "i";
ram[31] = "n";
ram[32] = " ";
ram[33] = "p";
ram[34] = "o";
ram[35] = "o";
ram[36] = "r";
ram[37] = " ";
ram[38] = "h";
ram[39] = "e";
ram[40] = "a";
ram[41] = "l";
ram[42] = "t";
ram[43] = "h";
ram[44] = ",";
ram[45] = " ";
ram[46] = "a";
ram[47] = "n";
ram[48] = "d";
ram[49] = " ";
ram[50] = "y";
ram[51] = "o";
ram[52] = "u";
ram[53] = " ";
ram[54] = "d";
ram[55] = "i";
ram[56] = "e";
ram[57] = " ";
ram[58] = "o";
ram[59] = "f";
ram[60] = " ";
ram[61] = "a";
ram[62] = " ";
ram[63] = "h";
ram[64] = "e";
ram[65] = "a";
ram[66] = "r";
ram[67] = "t";
ram[68] = " ";
ram[69] = "a";
ram[70] = "t";
ram[71] = "t";
ram[72] = "a";
ram[73] = "c";
ram[74] = "k";
ram[75] = ".";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
52 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "t";
ram[5] = "r";
ram[6] = "e";
ram[7] = "a";
ram[8] = "s";
ram[9] = "u";
ram[10] = "r";
ram[11] = "y";
ram[12] = " ";
ram[13] = "i";
ram[14] = "s";
ram[15] = " ";
ram[16] = "e";
ram[17] = "m";
ram[18] = "p";
ram[19] = "t";
ram[20] = "y";
ram[21] = ",";
ram[22] = " ";
ram[23] = "a";
ram[24] = "n";
ram[25] = "d";
ram[26] = " ";
ram[27] = "t";
ram[28] = "h";
ram[29] = "e";
ram[30] = " ";
ram[31] = "k";
ram[32] = "i";
ram[33] = "n";
ram[34] = "g";
ram[35] = "d";
ram[36] = "o";
ram[37] = "m";
ram[38] = " ";
ram[39] = "i";
ram[40] = "s";
ram[41] = " ";
ram[42] = "i";
ram[43] = "n";
ram[44] = " ";
ram[45] = "s";
ram[46] = "h";
ram[47] = "a";
ram[48] = "m";
ram[49] = "b";
ram[50] = "l";
ram[51] = "e";
ram[52] = "s";
ram[53] = ".";
ram[54] = " ";
ram[55] = "Y";
ram[56] = "o";
ram[57] = "u";
ram[58] = " ";
ram[59] = "d";
ram[60] = "i";
ram[61] = "e";
ram[62] = " ";
ram[63] = "o";
ram[64] = "f";
ram[65] = " ";
ram[66] = "m";
ram[67] = "a";
ram[68] = "l";
ram[69] = "n";
ram[70] = "u";
ram[71] = "t";
ram[72] = "r";
ram[73] = "i";
ram[74] = "t";
ram[75] = "i";
ram[76] = "o";
ram[77] = "n";
ram[78] = ".";
ram[79] = " ";
end
53 : begin
ram[0] = "Y";
ram[1] = "o";
ram[2] = "u";
ram[3] = "r";
ram[4] = " ";
ram[5] = "p";
ram[6] = "e";
ram[7] = "o";
ram[8] = "p";
ram[9] = "l";
ram[10] = "e";
ram[11] = " ";
ram[12] = "a";
ram[13] = "r";
ram[14] = "e";
ram[15] = " ";
ram[16] = "s";
ram[17] = "t";
ram[18] = "r";
ram[19] = "o";
ram[20] = "n";
ram[21] = "g";
ram[22] = " ";
ram[23] = "a";
ram[24] = "n";
ram[25] = "d";
ram[26] = " ";
ram[27] = "h";
ram[28] = "e";
ram[29] = "a";
ram[30] = "l";
ram[31] = "t";
ram[32] = "h";
ram[33] = "y";
ram[34] = ".";
ram[35] = " ";
ram[36] = "T";
ram[37] = "h";
ram[38] = "e";
ram[39] = "y";
ram[40] = " ";
ram[41] = "d";
ram[42] = "e";
ram[43] = "c";
ram[44] = "i";
ram[45] = "d";
ram[46] = "e";
ram[47] = " ";
ram[48] = "t";
ram[49] = "o";
ram[50] = " ";
ram[51] = "e";
ram[52] = "s";
ram[53] = "t";
ram[54] = "a";
ram[55] = "b";
ram[56] = "l";
ram[57] = "i";
ram[58] = "s";
ram[59] = "h";
ram[60] = " ";
ram[61] = "a";
ram[62] = " ";
ram[63] = "d";
ram[64] = "e";
ram[65] = "m";
ram[66] = "o";
ram[67] = "c";
ram[68] = "r";
ram[69] = "a";
ram[70] = "c";
ram[71] = "y";
ram[72] = ".";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
54 : begin
ram[0] = "Y";
ram[1] = "o";
ram[2] = "u";
ram[3] = " ";
ram[4] = "h";
ram[5] = "a";
ram[6] = "v";
ram[7] = "e";
ram[8] = " ";
ram[9] = "n";
ram[10] = "e";
ram[11] = "g";
ram[12] = "l";
ram[13] = "e";
ram[14] = "c";
ram[15] = "t";
ram[16] = "e";
ram[17] = "d";
ram[18] = " ";
ram[19] = "y";
ram[20] = "o";
ram[21] = "u";
ram[22] = "r";
ram[23] = " ";
ram[24] = "p";
ram[25] = "e";
ram[26] = "o";
ram[27] = "p";
ram[28] = "l";
ram[29] = "e";
ram[30] = ".";
ram[31] = " ";
ram[32] = "T";
ram[33] = "h";
ram[34] = "e";
ram[35] = "y";
ram[36] = " ";
ram[37] = "b";
ram[38] = "r";
ram[39] = "e";
ram[40] = "a";
ram[41] = "k";
ram[42] = " ";
ram[43] = "i";
ram[44] = "n";
ram[45] = "t";
ram[46] = "o";
ram[47] = " ";
ram[48] = "t";
ram[49] = "h";
ram[50] = "e";
ram[51] = " ";
ram[52] = "p";
ram[53] = "a";
ram[54] = "l";
ram[55] = "a";
ram[56] = "c";
ram[57] = "e";
ram[58] = " ";
ram[59] = "a";
ram[60] = "n";
ram[61] = "d";
ram[62] = " ";
ram[63] = "m";
ram[64] = "a";
ram[65] = "i";
ram[66] = "m";
ram[67] = " ";
ram[68] = "y";
ram[69] = "o";
ram[70] = "u";
ram[71] = ".";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
55 : begin
ram[0] = "Y";
ram[1] = "o";
ram[2] = "u";
ram[3] = "r";
ram[4] = " ";
ram[5] = "g";
ram[6] = "e";
ram[7] = "n";
ram[8] = "e";
ram[9] = "r";
ram[10] = "a";
ram[11] = "l";
ram[12] = "s";
ram[13] = " ";
ram[14] = "g";
ram[15] = "r";
ram[16] = "o";
ram[17] = "w";
ram[18] = " ";
ram[19] = "t";
ram[20] = "o";
ram[21] = "o";
ram[22] = " ";
ram[23] = "p";
ram[24] = "o";
ram[25] = "w";
ram[26] = "e";
ram[27] = "r";
ram[28] = "f";
ram[29] = "u";
ram[30] = "l";
ram[31] = ",";
ram[32] = " ";
ram[33] = "a";
ram[34] = "n";
ram[35] = "d";
ram[36] = " ";
ram[37] = "l";
ram[38] = "e";
ram[39] = "a";
ram[40] = "d";
ram[41] = " ";
ram[42] = "a";
ram[43] = " ";
ram[44] = "c";
ram[45] = "o";
ram[46] = "u";
ram[47] = "p";
ram[48] = ".";
ram[49] = " ";
ram[50] = "Y";
ram[51] = "o";
ram[52] = "u";
ram[53] = " ";
ram[54] = "a";
ram[55] = "r";
ram[56] = "e";
ram[57] = " ";
ram[58] = "k";
ram[59] = "i";
ram[60] = "l";
ram[61] = "l";
ram[62] = "e";
ram[63] = "d";
ram[64] = " ";
ram[65] = "i";
ram[66] = "n";
ram[67] = " ";
ram[68] = "t";
ram[69] = "h";
ram[70] = "e";
ram[71] = " ";
ram[72] = "c";
ram[73] = "h";
ram[74] = "a";
ram[75] = "o";
ram[76] = "s";
ram[77] = ".";
ram[78] = " ";
ram[79] = " ";
end
56 : begin
ram[0] = "Y";
ram[1] = "o";
ram[2] = "u";
ram[3] = " ";
ram[4] = "a";
ram[5] = "r";
ram[6] = "e";
ram[7] = " ";
ram[8] = "v";
ram[9] = "u";
ram[10] = "l";
ram[11] = "n";
ram[12] = "e";
ram[13] = "r";
ram[14] = "a";
ram[15] = "b";
ram[16] = "l";
ram[17] = "e";
ram[18] = " ";
ram[19] = "w";
ram[20] = "i";
ram[21] = "t";
ram[22] = "h";
ram[23] = "o";
ram[24] = "u";
ram[25] = "t";
ram[26] = " ";
ram[27] = "a";
ram[28] = "n";
ram[29] = " ";
ram[30] = "a";
ram[31] = "r";
ram[32] = "m";
ram[33] = "y";
ram[34] = ".";
ram[35] = " ";
ram[36] = "N";
ram[37] = "e";
ram[38] = "i";
ram[39] = "g";
ram[40] = "h";
ram[41] = "b";
ram[42] = "o";
ram[43] = "u";
ram[44] = "r";
ram[45] = "i";
ram[46] = "n";
ram[47] = "g";
ram[48] = " ";
ram[49] = "n";
ram[50] = "a";
ram[51] = "t";
ram[52] = "i";
ram[53] = "o";
ram[54] = "n";
ram[55] = "s";
ram[56] = " ";
ram[57] = "a";
ram[58] = "t";
ram[59] = "t";
ram[60] = "a";
ram[61] = "c";
ram[62] = "k";
ram[63] = " ";
ram[64] = "a";
ram[65] = "n";
ram[66] = "d";
ram[67] = " ";
ram[68] = "k";
ram[69] = "i";
ram[70] = "l";
ram[71] = "l";
ram[72] = " ";
ram[73] = "y";
ram[74] = "o";
ram[75] = "u";
ram[76] = ".";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
57 : begin
ram[0] = "T";
ram[1] = "h";
ram[2] = "e";
ram[3] = " ";
ram[4] = "c";
ram[5] = "h";
ram[6] = "u";
ram[7] = "r";
ram[8] = "c";
ram[9] = "h";
ram[10] = " ";
ram[11] = "g";
ram[12] = "r";
ram[13] = "o";
ram[14] = "w";
ram[15] = "s";
ram[16] = " ";
ram[17] = "t";
ram[18] = "o";
ram[19] = "o";
ram[20] = " ";
ram[21] = "p";
ram[22] = "o";
ram[23] = "w";
ram[24] = "e";
ram[25] = "r";
ram[26] = "f";
ram[27] = "u";
ram[28] = "l";
ram[29] = ",";
ram[30] = " ";
ram[31] = "a";
ram[32] = "n";
ram[33] = "d";
ram[34] = " ";
ram[35] = "o";
ram[36] = "v";
ram[37] = "e";
ram[38] = "r";
ram[39] = "t";
ram[40] = "h";
ram[41] = "r";
ram[42] = "o";
ram[43] = "w";
ram[44] = "s";
ram[45] = " ";
ram[46] = "t";
ram[47] = "h";
ram[48] = "e";
ram[49] = " ";
ram[50] = "m";
ram[51] = "o";
ram[52] = "n";
ram[53] = "a";
ram[54] = "r";
ram[55] = "c";
ram[56] = "h";
ram[57] = "y";
ram[58] = ".";
ram[59] = " ";
ram[60] = "Y";
ram[61] = "o";
ram[62] = "u";
ram[63] = " ";
ram[64] = "a";
ram[65] = "r";
ram[66] = "e";
ram[67] = " ";
ram[68] = "e";
ram[69] = "x";
ram[70] = "e";
ram[71] = "c";
ram[72] = "u";
ram[73] = "t";
ram[74] = "e";
ram[75] = "d";
ram[76] = ".";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
58 : begin
ram[0] = "Y";
ram[1] = "o";
ram[2] = "u";
ram[3] = " ";
ram[4] = "h";
ram[5] = "a";
ram[6] = "v";
ram[7] = "e";
ram[8] = " ";
ram[9] = "a";
ram[10] = "l";
ram[11] = "l";
ram[12] = "o";
ram[13] = "w";
ram[14] = "e";
ram[15] = "d";
ram[16] = " ";
ram[17] = "s";
ram[18] = "i";
ram[19] = "n";
ram[20] = " ";
ram[21] = "t";
ram[22] = "o";
ram[23] = " ";
ram[24] = "s";
ram[25] = "p";
ram[26] = "r";
ram[27] = "e";
ram[28] = "a";
ram[29] = "d";
ram[30] = " ";
ram[31] = "a";
ram[32] = "c";
ram[33] = "r";
ram[34] = "o";
ram[35] = "s";
ram[36] = "s";
ram[37] = " ";
ram[38] = "t";
ram[39] = "h";
ram[40] = "i";
ram[41] = "s";
ram[42] = " ";
ram[43] = "k";
ram[44] = "i";
ram[45] = "n";
ram[46] = "g";
ram[47] = "d";
ram[48] = "o";
ram[49] = "m";
ram[50] = ",";
ram[51] = " ";
ram[52] = "a";
ram[53] = "n";
ram[54] = "d";
ram[55] = " ";
ram[56] = "a";
ram[57] = "r";
ram[58] = "e";
ram[59] = " ";
ram[60] = "k";
ram[61] = "i";
ram[62] = "l";
ram[63] = "l";
ram[64] = "e";
ram[65] = "d";
ram[66] = " ";
ram[67] = "b";
ram[68] = "y";
ram[69] = " ";
ram[70] = "c";
ram[71] = "u";
ram[72] = "l";
ram[73] = "t";
ram[74] = "i";
ram[75] = "s";
ram[76] = "t";
ram[77] = "s";
ram[78] = ".";
ram[79] = " ";
end
59 : begin
ram[0] = "Y";
ram[1] = "o";
ram[2] = "u";
ram[3] = "r";
ram[4] = " ";
ram[5] = "M";
ram[6] = "a";
ram[7] = "j";
ram[8] = "e";
ram[9] = "s";
ram[10] = "t";
ram[11] = "y";
ram[12] = ",";
ram[13] = " ";
ram[14] = "w";
ram[15] = "a";
ram[16] = "k";
ram[17] = "e";
ram[18] = " ";
ram[19] = "u";
ram[20] = "p";
ram[21] = "!";
ram[22] = " ";
ram[23] = "Y";
ram[24] = "o";
ram[25] = "u";
ram[26] = "r";
ram[27] = " ";
ram[28] = "l";
ram[29] = "o";
ram[30] = "y";
ram[31] = "a";
ram[32] = "l";
ram[33] = " ";
ram[34] = "s";
ram[35] = "u";
ram[36] = "b";
ram[37] = "j";
ram[38] = "e";
ram[39] = "c";
ram[40] = "t";
ram[41] = "s";
ram[42] = " ";
ram[43] = "n";
ram[44] = "e";
ram[45] = "e";
ram[46] = "d";
ram[47] = " ";
ram[48] = "g";
ram[49] = "u";
ram[50] = "i";
ram[51] = "d";
ram[52] = "a";
ram[53] = "n";
ram[54] = "c";
ram[55] = "e";
ram[56] = " ";
ram[57] = "o";
ram[58] = "n";
ram[59] = " ";
ram[60] = "s";
ram[61] = "t";
ram[62] = "a";
ram[63] = "t";
ram[64] = "e";
ram[65] = "l";
ram[66] = "y";
ram[67] = " ";
ram[68] = "a";
ram[69] = "f";
ram[70] = "f";
ram[71] = "a";
ram[72] = "i";
ram[73] = "r";
ram[74] = "s";
ram[75] = ".";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
60 : begin
ram[0] = "I";
ram[1] = " ";
ram[2] = "A";
ram[3] = "M";
ram[4] = " ";
ram[5] = "A";
ram[6] = " ";
ram[7] = "F";
ram[8] = "I";
ram[9] = "L";
ram[10] = "E";
ram[11] = " ";
ram[12] = "A";
ram[13] = "N";
ram[14] = "D";
ram[15] = " ";
ram[16] = "Y";
ram[17] = "O";
ram[18] = "U";
ram[19] = " ";
ram[20] = "P";
ram[21] = "U";
ram[22] = "T";
ram[23] = " ";
ram[24] = "D";
ram[25] = "O";
ram[26] = "C";
ram[27] = "U";
ram[28] = "M";
ram[29] = "E";
ram[30] = "N";
ram[31] = "T";
ram[32] = "S";
ram[33] = " ";
ram[34] = "I";
ram[35] = "N";
ram[36] = " ";
ram[37] = "M";
ram[38] = "E";
ram[39] = ".";
ram[40] = "I";
ram[41] = " ";
ram[42] = "A";
ram[43] = "M";
ram[44] = " ";
ram[45] = "A";
ram[46] = " ";
ram[47] = "F";
ram[48] = "I";
ram[49] = "L";
ram[50] = "E";
ram[51] = " ";
ram[52] = "A";
ram[53] = "N";
ram[54] = "D";
ram[55] = " ";
ram[56] = "Y";
ram[57] = "O";
ram[58] = "U";
ram[59] = " ";
ram[60] = "P";
ram[61] = "U";
ram[62] = "T";
ram[63] = " ";
ram[64] = "D";
ram[65] = "O";
ram[66] = "C";
ram[67] = "U";
ram[68] = "M";
ram[69] = "E";
ram[70] = "N";
ram[71] = "T";
ram[72] = "S";
ram[73] = " ";
ram[74] = "I";
ram[75] = "N";
ram[76] = " ";
ram[77] = "M";
ram[78] = "E";
ram[79] = ".";
end
61 : begin
ram[0] = "Y";
ram[1] = "o";
ram[2] = "u";
ram[3] = " ";
ram[4] = "h";
ram[5] = "a";
ram[6] = "v";
ram[7] = "e";
ram[8] = " ";
ram[9] = "r";
ram[10] = "u";
ram[11] = "l";
ram[12] = "e";
ram[13] = "d";
ram[14] = " ";
ram[15] = "w";
ram[16] = "e";
ram[17] = "l";
ram[18] = "l";
ram[19] = " ";
ram[20] = "f";
ram[21] = "o";
ram[22] = "r";
ram[23] = " ";
ram[24] = "5";
ram[25] = "0";
ram[26] = " ";
ram[27] = "y";
ram[28] = "e";
ram[29] = "a";
ram[30] = "r";
ram[31] = "s";
ram[32] = ".";
ram[33] = " ";
ram[34] = "Y";
ram[35] = "o";
ram[36] = "u";
ram[37] = " ";
ram[38] = "p";
ram[39] = "a";
ram[40] = "s";
ram[41] = "s";
ram[42] = " ";
ram[43] = "a";
ram[44] = "w";
ram[45] = "a";
ram[46] = "y";
ram[47] = " ";
ram[48] = "p";
ram[49] = "e";
ram[50] = "a";
ram[51] = "c";
ram[52] = "e";
ram[53] = "f";
ram[54] = "u";
ram[55] = "l";
ram[56] = "l";
ram[57] = "y";
ram[58] = ",";
ram[59] = " ";
ram[60] = "l";
ram[61] = "o";
ram[62] = "v";
ram[63] = "e";
ram[64] = "d";
ram[65] = " ";
ram[66] = "b";
ram[67] = "y";
ram[68] = " ";
ram[69] = "a";
ram[70] = "l";
ram[71] = "l";
ram[72] = ".";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end
62 : begin
ram[0] = "S";
ram[1] = "e";
ram[2] = "l";
ram[3] = "e";
ram[4] = "c";
ram[5] = "t";
ram[6] = " ";
ram[7] = "y";
ram[8] = "o";
ram[9] = "u";
ram[10] = "r";
ram[11] = " ";
ram[12] = "d";
ram[13] = "i";
ram[14] = "f";
ram[15] = "f";
ram[16] = "i";
ram[17] = "c";
ram[18] = "u";
ram[19] = "l";
ram[20] = "t";
ram[21] = "y";
ram[22] = " ";
ram[23] = "m";
ram[24] = "y";
ram[25] = " ";
ram[26] = "l";
ram[27] = "i";
ram[28] = "e";
ram[29] = "g";
ram[30] = "e";
ram[31] = ".";
ram[32] = " ";
ram[33] = " ";
ram[34] = " ";
ram[35] = " ";
ram[36] = " ";
ram[37] = " ";
ram[38] = " ";
ram[39] = " ";
ram[40] = " ";
ram[41] = " ";
ram[42] = "N";
ram[43] = "O";
ram[44] = "R";
ram[45] = "M";
ram[46] = "A";
ram[47] = "L";
ram[48] = " ";
ram[49] = " ";
ram[50] = " ";
ram[51] = " ";
ram[52] = " ";
ram[53] = " ";
ram[54] = " ";
ram[55] = " ";
ram[56] = " ";
ram[57] = " ";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = "A";
ram[72] = "N";
ram[73] = "A";
ram[74] = "R";
ram[75] = "C";
ram[76] = "H";
ram[77] = "Y";
ram[78] = " ";
ram[79] = " ";
end
63 : begin
ram[0] = "W";
ram[1] = "e";
ram[2] = "l";
ram[3] = "c";
ram[4] = "o";
ram[5] = "m";
ram[6] = "e";
ram[7] = ",";
ram[8] = " ";
ram[9] = "Y";
ram[10] = "o";
ram[11] = "u";
ram[12] = "r";
ram[13] = " ";
ram[14] = "M";
ram[15] = "a";
ram[16] = "j";
ram[17] = "e";
ram[18] = "s";
ram[19] = "t";
ram[20] = "y";
ram[21] = "!";
ram[22] = " ";
ram[23] = "P";
ram[24] = "r";
ram[25] = "e";
ram[26] = "s";
ram[27] = "s";
ram[28] = " ";
ram[29] = "a";
ram[30] = "n";
ram[31] = "y";
ram[32] = " ";
ram[33] = "k";
ram[34] = "e";
ram[35] = "y";
ram[36] = " ";
ram[37] = "t";
ram[38] = "o";
ram[39] = " ";
ram[40] = "s";
ram[41] = "t";
ram[42] = "a";
ram[43] = "r";
ram[44] = "t";
ram[45] = ".";
ram[46] = " ";
ram[47] = " ";
ram[48] = " ";
ram[49] = " ";
ram[50] = " ";
ram[51] = " ";
ram[52] = " ";
ram[53] = " ";
ram[54] = " ";
ram[55] = " ";
ram[56] = " ";
ram[57] = " ";
ram[58] = " ";
ram[59] = " ";
ram[60] = " ";
ram[61] = " ";
ram[62] = " ";
ram[63] = " ";
ram[64] = " ";
ram[65] = " ";
ram[66] = " ";
ram[67] = " ";
ram[68] = " ";
ram[69] = " ";
ram[70] = " ";
ram[71] = " ";
ram[72] = " ";
ram[73] = " ";
ram[74] = " ";
ram[75] = " ";
ram[76] = " ";
ram[77] = " ";
ram[78] = " ";
ram[79] = " ";
end

endcase

end
  
  always @(posedge clk) begin
    read_data <= ram[address];         // read the entry
    
    if (write_en)                      // if we need to write
      ram[address] <= write_data;      // update that value
  end
  
endmodule